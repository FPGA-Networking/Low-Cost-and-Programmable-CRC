// **************************************************************
// COPYRIGHT(c)2015, Xidian University
// All rights reserved.
//
// IP LIB INDEX :  
// IP Name      :      
// File name    : 
// Module name  : 
// Full name    :  
//
// Author       : Liu-Huan 
// Email        : assasin9997@163.com 
// Data         : 
// Version      : V 1.0 
// 
// Abstract     : 
// Called by    :  
// 
// Modification history
// -----------------------------------------------------------------
// 
// 
//
// *****************************************************************

// *******************
// TIMESCALE
// ******************* 
`timescale 1ns/1ps 

// *******************
// INFORMATION
// *******************


//*******************
//DEFINE(s)
//*******************
//`define UDLY 1    //Unit delay, for non-blocking assignments in sequential logic



//*******************
//DEFINE MODULE PORT
//*******************
module  go_back_top  

# ( parameter   
                SEG_NUM              = 0 ,
                BUS_WIDTH            = 0 ,
                BUS_WIDTH_MULTI_6    = 0 ,
                MOD_WIDTH            = 0 ,
                CMP_LAYER            = 0 ,      // C_XOR之前计算的层数，包含第一层
                GO_BACK_STAGE        = 0 ,
                LUT_NUM_LAYER_1      = 0 ,
                LUT_NUM_LAYER_2      = 0 ,
                LUT_NUM_LAYER_3      = 0 ,
                LUT_NUM_LAYER_4      = 0 ,
                LUT_NUM_LAYER_5      = 0 ,
                LUT_NUM_LAYER_6      = 0 ,
                LUT_NUM_LAYER_7      = 0 ,
                LUT_NUM_LAYER_8      = 0 ,                
                LUT_OUT_NUM_LAYER_1  = 0 ,
                LUT_OUT_NUM_LAYER_2  = 0 ,
                LUT_OUT_NUM_LAYER_3  = 0 ,
                LUT_OUT_NUM_LAYER_4  = 0 ,
                LUT_OUT_NUM_LAYER_5  = 0 ,
                LUT_OUT_NUM_LAYER_6  = 0 ,
                LUT_OUT_NUM_LAYER_7  = 0 ,
                LUT_OUT_NUM_LAYER_8  = 0 ,
                PKT_NUM              = 0    
        )
  (     
            input                           clk  ,
            input                           rst  ,
            input  [SEG_NUM-1:0]            seg_sop        ,
            input  [SEG_NUM-1:0]            seg_eop        ,
            input  [SEG_NUM-1:0]            seg_dval       ,
            input  [SEG_NUM*4-1:0]          seg_packet_num ,
            input  [SEG_NUM*12-1:0]         seg_zero_num   ,
            input  [SEG_NUM*BUS_WIDTH-1:0]  seg_dout       , 

            output   [PKT_NUM-1:0]            crc_en  ,
            output   [32*PKT_NUM-1:0]         crc 


              ) ;



parameter  [0:SEG_NUM*LUT_NUM_LAYER_1*64*16-1] D_LUT_POLY = {

64'b1010101010101010101010101010101001010101010101011010101010101010,
64'b0011001100110011110011001100110001010101101010100101010110101010,
64'b0101101001011010010110100101101000001111111100000000111111110000,
64'b1100110011001100110011001100110000001111000011111111000011110000,
64'b1111111111111111000000000000000011000011110000110011110000111100,
64'b0110011010011001100110010110011000110011001100111100110011001100,
64'b0110100101101001100101101001011001011010010110100101101001011010,
64'b1111000011110000111100001111000001011010010110100101101001011010,
64'b1111111111111111000000000000000011111111111111110000000000000000,
64'b1010010101011010101001010101101011000011001111001100001100111100,
64'b1010101001010101010101011010101011001100110011001100110011001100,
64'b0101010110101010010101011010101000111100001111000011110000111100,
64'b1001100101100110100110010110011000000000000000000000000000000000,
64'b0110011001100110011001100110011011001100110011001100110011001100,
64'b1100001111000011001111000011110010011001100110010110011001100110,
64'b1100001100111100110000110011110000000000111111111111111100000000,
64'b0011110000111100001111000011110011111111000000001111111100000000,
64'b1111111111111111000000000000000010100101010110101010010101011010,
64'b0000111111110000000011111111000001011010010110100101101001011010,
64'b0000000011111111111111110000000010011001011001101001100101100110,
64'b1010010101011010101001010101101000110011110011000011001111001100,
64'b1111111111111111000000000000000000000000000000000000000000000000,
64'b1100001111000011001111000011110001011010101001011010010101011010,
64'b1001100101100110100110010110011011110000111100001111000011110000,
64'b1100110000110011001100111100110000001111111100000000111111110000,
64'b1010010101011010101001010101101000000000000000000000000000000000,
64'b1001011010010110100101101001011011110000111100001111000011110000,
64'b0011110011000011110000110011110000111100001111000011110000111100,
64'b0000000011111111111111110000000001010101010101011010101010101010,
64'b1100001100111100110000110011110001010101010101011010101010101010,
64'b1111111111111111000000000000000011001100001100110011001111001100,
64'b1100110011001100110011001100110000110011110011000011001111001100,
64'b1001011010010110100101101001011011000011110000110011110000111100,
64'b1001011001101001011010011001011000001111000011111111000011110000,
64'b1111111111111111000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000011001100001100110011001111001100,
64'b1100001100111100110000110011110001010101101010100101010110101010,
64'b0101101010100101101001010101101000000000111111111111111100000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1100001100111100110000110011110011111111000000001111111100000000,
64'b1111000000001111000011111111000000001111111100000000111111110000,
64'b0101010101010101101010101010101011001100110011001100110011001100,
64'b0101101010100101101001010101101001100110011001100110011001100110,
64'b0000000000000000000000000000000010100101101001010101101001011010,
64'b0101101001011010010110100101101010100101101001010101101001011010,
64'b1100001100111100110000110011110000001111111100000000111111110000,
64'b0011110011000011110000110011110001010101101010100101010110101010,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b1010101010101010101010101010101000001111000011111111000011110000,
64'b1111000000001111000011111111000010011001100110010110011001100110,
64'b1100110000110011001100111100110011111111111111110000000000000000,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b0101101010100101101001010101101011111111111111110000000000000000,
64'b0011001111001100001100111100110000000000111111111111111100000000,
64'b0011110000111100001111000011110011110000111100001111000011110000,
64'b1010101001010101010101011010101000111100001111000011110000111100,
64'b0101010101010101101010101010101000110011110011000011001111001100,
64'b0101010101010101101010101010101010011001011001101001100101100110,
64'b1001100101100110100110010110011010101010010101010101010110101010,
64'b0000000011111111111111110000000000110011001100111100110011001100,
64'b1001100110011001011001100110011011001100110011001100110011001100,
64'b0110100110010110011010011001011011111111000000001111111100000000,
64'b1010101010101010101010101010101010010110100101101001011010010110,
64'b1111000000001111000011111111000010101010101010101010101010101010,
64'b1111111100000000111111110000000001100110011001100110011001100110,
64'b0110011010011001100110010110011000000000000000000000000000000000,
64'b1001011010010110100101101001011001010101010101011010101010101010,
64'b0101010110101010010101011010101001010101101010100101010110101010,
64'b1111111111111111000000000000000000001111111100000000111111110000,
64'b1001100110011001011001100110011000001111000011111111000011110000,
64'b0000000011111111111111110000000011000011110000110011110000111100,
64'b0000000000000000000000000000000000110011001100111100110011001100,
64'b0000111100001111111100001111000001011010010110100101101001011010,
64'b0110100101101001100101101001011001011010010110100101101001011010,
64'b0011001100110011110011001100110011111111111111110000000000000000,
64'b0110011010011001100110010110011011000011001111001100001100111100,
64'b0101010101010101101010101010101011001100110011001100110011001100,
64'b0011001111001100001100111100110000111100001111000011110000111100,
64'b1100001111000011001111000011110010101010101010101010101010101010,
64'b0110100110010110011010011001011011111111111111110000000000000000,
64'b0011001100110011110011001100110011000011110000110011110000111100,
64'b0000000000000000000000000000000011001100001100110011001111001100,
64'b1001011010010110100101101001011000000000111111111111111100000000,
64'b0101010101010101101010101010101011000011110000110011110000111100,
64'b1010101010101010101010101010101000110011001100111100110011001100,
64'b1111111100000000111111110000000001101001100101100110100110010110,
64'b0110100110010110011010011001011011001100001100110011001111001100,
64'b0101101001011010010110100101101010100101010110101010010101011010,
64'b0110100101101001100101101001011011110000111100001111000011110000,
64'b0110011001100110011001100110011010100101010110101010010101011010,
64'b0101101001011010010110100101101010010110100101101001011010010110,
64'b1010010101011010101001010101101001100110011001100110011001100110,
64'b1010010101011010101001010101101000110011001100111100110011001100,
64'b1010101010101010101010101010101011111111000000001111111100000000,
64'b0110011001100110011001100110011001101001011010011001011010010110,
64'b0011110011000011110000110011110010101010101010101010101010101010,
64'b1010101001010101010101011010101011000011110000110011110000111100,
64'b0000111100001111111100001111000000110011001100111100110011001100,
64'b0000111100001111111100001111000001100110100110011001100101100110,
64'b1100001100111100110000110011110011110000111100001111000011110000,
64'b1001011010010110100101101001011011000011110000110011110000111100,
64'b0110100101101001100101101001011001010101010101011010101010101010,
64'b1100001100111100110000110011110010011001100110010110011001100110,
64'b1010101010101010101010101010101001011010010110100101101001011010,
64'b0110011010011001100110010110011000111100001111000011110000111100,
64'b1111111100000000111111110000000011110000111100001111000011110000,
64'b1001011010010110100101101001011001010101010101011010101010101010,
64'b1111000011110000111100001111000011000011001111001100001100111100,
64'b0000111111110000000011111111000001100110011001100110011001100110,
64'b1111111100000000111111110000000000001111111100000000111111110000,
64'b0011110011000011110000110011110001011010010110100101101001011010,
64'b1010010101011010101001010101101001101001011010011001011010010110,
64'b1010010101011010101001010101101001010101101010100101010110101010,
64'b0110011001100110011001100110011000001111111100000000111111110000,
64'b0110100101101001100101101001011001100110011001100110011001100110,
64'b0000111100001111111100001111000010010110100101101001011010010110,
64'b0101010110101010010101011010101010011001011001101001100101100110,
64'b1100001111000011001111000011110000001111111100000000111111110000,
64'b0101010101010101101010101010101011111111000000001111111100000000,
64'b1100001100111100110000110011110011001100110011001100110011001100,
64'b1111111100000000111111110000000001011010101001011010010101011010,
64'b0000000011111111111111110000000000111100001111000011110000111100,
64'b1111111111111111000000000000000000000000111111111111111100000000,
64'b1111000000001111000011111111000000110011110011000011001111001100,
64'b0110011010011001100110010110011011000011001111001100001100111100,
64'b1100110000110011001100111100110010011001100110010110011001100110,
64'b0011110000111100001111000011110000000000111111111111111100000000,
64'b1100001100111100110000110011110000111100001111000011110000111100,
64'b0101010110101010010101011010101011000011001111001100001100111100,
64'b0110011001100110011001100110011000111100001111000011110000111100,
64'b1010010101011010101001010101101010101010010101010101010110101010,
64'b0101010101010101101010101010101011001100110011001100110011001100,
64'b0000000011111111111111110000000010101010101010101010101010101010,
64'b0011001100110011110011001100110000000000111111111111111100000000,
64'b0000000000000000000000000000000001011010101001011010010101011010,
64'b1100110000110011001100111100110010011001011001101001100101100110,
64'b1100001100111100110000110011110011001100110011001100110011001100,
64'b1001100110011001011001100110011000000000111111111111111100000000,
64'b0101101001011010010110100101101011000011110000110011110000111100,
64'b0000000000000000000000000000000011110000000011110000111111110000,
64'b0101101001011010010110100101101000001111000011111111000011110000,
64'b0110011010011001100110010110011010100101101001010101101001011010,
64'b1010010101011010101001010101101010010110100101101001011010010110,
64'b0110011010011001100110010110011000110011001100111100110011001100,
64'b1111111111111111000000000000000001011010010110100101101001011010,
64'b0000111100001111111100001111000011001100110011001100110011001100,
64'b1001011010010110100101101001011011111111111111110000000000000000,
64'b0101010101010101101010101010101001100110100110011001100101100110,
64'b0110100110010110011010011001011001101001011010011001011010010110,
64'b0011001111001100001100111100110011110000111100001111000011110000,
64'b1100110011001100110011001100110011111111111111110000000000000000,
64'b0110011010011001100110010110011010100101010110101010010101011010,
64'b1010010101011010101001010101101010101010010101010101010110101010,
64'b1001100110011001011001100110011001010101101010100101010110101010,
64'b1001011001101001011010011001011010011001011001101001100101100110,
64'b0000000000000000000000000000000001101001100101100110100110010110,
64'b0110100101101001100101101001011011110000111100001111000011110000,
64'b1001100110011001011001100110011010011001011001101001100101100110,
64'b0000111111110000000011111111000011110000111100001111000011110000,
64'b1010010101011010101001010101101000000000000000000000000000000000,
64'b0011001100110011110011001100110001101001011010011001011010010110,
64'b1111000011110000111100001111000001101001100101100110100110010110,
64'b0110011001100110011001100110011001010101101010100101010110101010,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0011110000111100001111000011110001100110100110011001100101100110,
64'b1100001111000011001111000011110000110011001100111100110011001100,
64'b1001011001101001011010011001011010011001100110010110011001100110,
64'b1100001111000011001111000011110011000011110000110011110000111100,
64'b0011001111001100001100111100110011000011001111001100001100111100,
64'b1100001100111100110000110011110011111111000000001111111100000000,
64'b1001011010010110100101101001011011000011110000110011110000111100,
64'b1010101001010101010101011010101011111111000000001111111100000000,
64'b1100110000110011001100111100110000000000000000000000000000000000,
64'b1111000011110000111100001111000011000011001111001100001100111100,
64'b0101010110101010010101011010101010010110011010010110100110010110,
64'b0011110000111100001111000011110000110011001100111100110011001100,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000111111110000000011111111000011000011110000110011110000111100,
64'b0000111111110000000011111111000001011010010110100101101001011010,
64'b1001011001101001011010011001011010010110100101101001011010010110,
64'b1010010101011010101001010101101010100101010110101010010101011010,
64'b0101101001011010010110100101101010100101010110101010010101011010,
64'b1111000000001111000011111111000011111111111111110000000000000000,
64'b1100001100111100110000110011110000001111111100000000111111110000,
64'b0011001100110011110011001100110001010101010101011010101010101010,
64'b1010010110100101010110100101101000000000000000000000000000000000,
64'b0101010110101010010101011010101011110000000011110000111111110000,
64'b0011001100110011110011001100110000111100110000111100001100111100,
64'b0000111111110000000011111111000001011010010110100101101001011010,
64'b0000000000000000000000000000000010101010101010101010101010101010,
64'b0000000011111111111111110000000000001111111100000000111111110000,
64'b0000000011111111111111110000000010011001011001101001100101100110,
64'b0011110011000011110000110011110011000011001111001100001100111100,
64'b0110011010011001100110010110011011001100001100110011001111001100,
64'b0011001111001100001100111100110000110011110011000011001111001100,
64'b0000000011111111111111110000000000000000000000000000000000000000,
64'b0101101010100101101001010101101010101010010101010101010110101010,
64'b1111000011110000111100001111000011001100110011001100110011001100,
64'b1001100101100110100110010110011010101010101010101010101010101010,
64'b1001100110011001011001100110011000000000111111111111111100000000,
64'b1111000011110000111100001111000001011010101001011010010101011010,
64'b1010101001010101010101011010101010011001011001101001100101100110,
64'b0000000000000000000000000000000011001100110011001100110011001100,
64'b1111111111111111000000000000000000000000111111111111111100000000,
64'b0101010101010101101010101010101011000011110000110011110000111100,
64'b0101101010100101101001010101101011110000000011110000111111110000,
64'b0110100101101001100101101001011000001111000011111111000011110000,
64'b0101101001011010010110100101101001011010010110100101101001011010,
64'b0011110011000011110000110011110000001111000011111111000011110000,
64'b0000000011111111111111110000000000000000000000000000000000000000,
64'b0000000000000000000000000000000011001100001100110011001111001100,
64'b0101101010100101101001010101101000000000111111111111111100000000,
64'b1001100101100110100110010110011010100101010110101010010101011010,
64'b0000000000000000000000000000000010010110100101101001011010010110,
64'b1001011001101001011010011001011001010101101010100101010110101010,
64'b1010010110100101010110100101101001100110100110011001100101100110,
64'b0101101001011010010110100101101001100110011001100110011001100110,
64'b1100001111000011001111000011110001101001100101100110100110010110,
64'b0101101010100101101001010101101011000011110000110011110000111100,
64'b0101010101010101101010101010101010010110100101101001011010010110,
64'b1100001100111100110000110011110001010101101010100101010110101010,
64'b0110011001100110011001100110011011111111000000001111111100000000,
64'b0101010110101010010101011010101010101010101010101010101010101010,
64'b1010101010101010101010101010101000001111000011111111000011110000,
64'b1001011010010110100101101001011001010101010101011010101010101010,
64'b1111000000001111000011111111000001100110100110011001100101100110,
64'b0000000000000000000000000000000011000011001111001100001100111100,
64'b1010101010101010101010101010101000110011001100111100110011001100,
64'b0011110011000011110000110011110011000011110000110011110000111100,
64'b1100001100111100110000110011110010010110100101101001011010010110,
64'b1100110000110011001100111100110000111100110000111100001100111100,
64'b0011110000111100001111000011110000001111111100000000111111110000,
64'b0011001100110011110011001100110001101001100101100110100110010110,
64'b0110011001100110011001100110011011001100110011001100110011001100,
64'b1010101001010101010101011010101011111111111111110000000000000000,
64'b0011001111001100001100111100110011001100110011001100110011001100,
64'b1100110011001100110011001100110011111111000000001111111100000000,
64'b1001100110011001011001100110011001100110011001100110011001100110,
64'b1001100110011001011001100110011001101001011010011001011010010110,
64'b1010101010101010101010101010101001011010101001011010010101011010,
64'b0101101010100101101001010101101011110000111100001111000011110000,
64'b0101010110101010010101011010101010100101010110101010010101011010,
64'b0000000011111111111111110000000001101001100101100110100110010110,
64'b1100110011001100110011001100110011110000000011110000111111110000,
64'b1111111111111111000000000000000010101010010101010101010110101010,
64'b1010010110100101010110100101101000111100110000111100001100111100,
64'b0101010110101010010101011010101011110000111100001111000011110000,
64'b0011001100110011110011001100110000000000000000000000000000000000,
64'b1010010110100101010110100101101001011010010110100101101001011010,
64'b1111000011110000111100001111000011111111111111110000000000000000,
64'b0011110000111100001111000011110000111100001111000011110000111100,
64'b1001011010010110100101101001011011000011001111001100001100111100,
64'b0110011001100110011001100110011001100110100110011001100101100110,
64'b1100110000110011001100111100110001010101101010100101010110101010,
64'b1001100110011001011001100110011011001100001100110011001111001100,
64'b1111111111111111000000000000000000111100110000111100001100111100,
64'b0101101001011010010110100101101000000000111111111111111100000000,
64'b0000000000000000000000000000000010011001100110010110011001100110,
64'b1001100101100110100110010110011001011010101001011010010101011010,
64'b0110011001100110011001100110011001010101101010100101010110101010,
64'b1100110000110011001100111100110000000000000000000000000000000000,
64'b1001100110011001011001100110011000110011110011000011001111001100,
64'b0101010110101010010101011010101000000000000000000000000000000000,
64'b0101010101010101101010101010101010100101010110101010010101011010,
64'b0101101001011010010110100101101011110000000011110000111111110000,
64'b0011110000111100001111000011110011000011110000110011110000111100,
64'b1001100101100110100110010110011010011001100110010110011001100110,
64'b0011001100110011110011001100110000001111000011111111000011110000,
64'b1111000011110000111100001111000001011010101001011010010101011010,
64'b0101101010100101101001010101101001010101010101011010101010101010,
64'b0101101010100101101001010101101010010110100101101001011010010110,
64'b1001011010010110100101101001011001100110100110011001100101100110,
64'b1111111100000000111111110000000001100110011001100110011001100110,
64'b1001100101100110100110010110011000000000000000000000000000000000,
64'b1001011001101001011010011001011000001111000011111111000011110000,
64'b1001100110011001011001100110011000000000000000000000000000000000,
64'b1001011001101001011010011001011011001100001100110011001111001100,
64'b0000000000000000000000000000000000000000111111111111111100000000,
64'b0000111111110000000011111111000010100101010110101010010101011010,
64'b0101010110101010010101011010101010010110100101101001011010010110,
64'b0101010101010101101010101010101001010101101010100101010110101010,
64'b0000111111110000000011111111000001100110100110011001100101100110,
64'b0000111111110000000011111111000001100110011001100110011001100110,
64'b0011110000111100001111000011110001101001100101100110100110010110,
64'b0011110011000011110000110011110011000011110000110011110000111100,
64'b1100001100111100110000110011110010010110100101101001011010010110,
64'b0110100101101001100101101001011000111100110000111100001100111100,
64'b0011110011000011110000110011110011111111111111110000000000000000,
64'b1001011010010110100101101001011010101010101010101010101010101010,
64'b1001011001101001011010011001011001010101101010100101010110101010,
64'b1010101010101010101010101010101011001100001100110011001111001100,
64'b0000000011111111111111110000000001100110100110011001100101100110,
64'b0011001100110011110011001100110001010101010101011010101010101010,
64'b1100110011001100110011001100110010010110100101101001011010010110,
64'b1010101001010101010101011010101010011001100110010110011001100110,
64'b0000000011111111111111110000000001010101010101011010101010101010,
64'b0000111111110000000011111111000001100110011001100110011001100110,
64'b1111000000001111000011111111000001011010101001011010010101011010,
64'b1010010101011010101001010101101010101010101010101010101010101010,
64'b1111111111111111000000000000000011001100110011001100110011001100,
64'b0101101001011010010110100101101010101010010101010101010110101010,
64'b0110100110010110011010011001011001100110011001100110011001100110,
64'b0110011001100110011001100110011001101001100101100110100110010110,
64'b1111111100000000111111110000000010010110011010010110100110010110,
64'b1111111111111111000000000000000001101001011010011001011010010110,
64'b1100110000110011001100111100110011110000000011110000111111110000,
64'b1111111111111111000000000000000011001100001100110011001111001100,
64'b0110100101101001100101101001011001100110011001100110011001100110,
64'b1001011010010110100101101001011010100101101001010101101001011010,
64'b1111000011110000111100001111000011001100001100110011001111001100,
64'b0101010110101010010101011010101010011001011001101001100101100110,
64'b0101101001011010010110100101101010100101010110101010010101011010,
64'b0011110011000011110000110011110011110000111100001111000011110000,
64'b1001100110011001011001100110011000110011001100111100110011001100,
64'b0011110011000011110000110011110010010110100101101001011010010110,
64'b0110011010011001100110010110011000111100110000111100001100111100,
64'b0110011010011001100110010110011000111100110000111100001100111100,
64'b0000000000000000000000000000000001101001100101100110100110010110,
64'b0011001111001100001100111100110010101010010101010101010110101010,
64'b0000111100001111111100001111000010100101101001010101101001011010,
64'b0011001111001100001100111100110010010110100101101001011010010110,
64'b1010101001010101010101011010101000110011110011000011001111001100,
64'b1010010110100101010110100101101010100101101001010101101001011010,
64'b0110011001100110011001100110011001101001011010011001011010010110,
64'b1111000011110000111100001111000000110011110011000011001111001100,
64'b0101101010100101101001010101101001010101101010100101010110101010,
64'b1001011010010110100101101001011011110000111100001111000011110000,
64'b0101101010100101101001010101101001101001100101100110100110010110,
64'b0110100101101001100101101001011011110000000011110000111111110000,
64'b0110100101101001100101101001011001011010101001011010010101011010,
64'b1010101010101010101010101010101010010110011010010110100110010110,
64'b0000111100001111111100001111000000110011001100111100110011001100,
64'b1111111100000000111111110000000010011001011001101001100101100110,
64'b1010010110100101010110100101101001101001100101100110100110010110,
64'b0011001100110011110011001100110000001111000011111111000011110000,
64'b1001100101100110100110010110011000110011110011000011001111001100,
64'b1001011010010110100101101001011001101001100101100110100110010110,
64'b1111111100000000111111110000000001011010010110100101101001011010,
64'b1111000011110000111100001111000000001111111100000000111111110000,
64'b0110100101101001100101101001011011111111111111110000000000000000,
64'b1100110000110011001100111100110000111100110000111100001100111100,
64'b0011001100110011110011001100110001011010010110100101101001011010,
64'b1111000011110000111100001111000011111111111111110000000000000000,
64'b0110011001100110011001100110011010010110011010010110100110010110,
64'b0110100101101001100101101001011011001100001100110011001111001100,
64'b1111000011110000111100001111000011001100110011001100110011001100,
64'b0110100110010110011010011001011001100110100110011001100101100110,
64'b1001100110011001011001100110011000111100110000111100001100111100,
64'b0011001111001100001100111100110011111111000000001111111100000000,
64'b1001011001101001011010011001011001101001100101100110100110010110,
64'b1100001100111100110000110011110011110000111100001111000011110000,
64'b0110100101101001100101101001011000000000111111111111111100000000,
64'b1100001111000011001111000011110000000000000000000000000000000000,
64'b1010010110100101010110100101101001011010101001011010010101011010,
64'b0000000011111111111111110000000010011001011001101001100101100110,
64'b1100110011001100110011001100110000000000000000000000000000000000,
64'b0011110000111100001111000011110010010110011010010110100110010110,
64'b0101010101010101101010101010101010100101101001010101101001011010,
64'b1111000000001111000011111111000001011010010110100101101001011010,
64'b0110011010011001100110010110011011000011110000110011110000111100,
64'b1111111111111111000000000000000001011010101001011010010101011010,
64'b1111111100000000111111110000000001010101010101011010101010101010,
64'b0110100110010110011010011001011000111100110000111100001100111100,
64'b0110011001100110011001100110011011111111000000001111111100000000,
64'b1111111111111111000000000000000001010101010101011010101010101010,
64'b1010010110100101010110100101101010101010101010101010101010101010,
64'b1001100101100110100110010110011011001100001100110011001111001100,
64'b0000111111110000000011111111000001101001011010011001011010010110,
64'b1100001100111100110000110011110000000000000000000000000000000000,
64'b0000111111110000000011111111000000111100110000111100001100111100,
64'b0101101010100101101001010101101010011001011001101001100101100110,
64'b0000111111110000000011111111000010011001011001101001100101100110,
64'b0011001100110011110011001100110000001111111100000000111111110000,
64'b0110100101101001100101101001011001100110100110011001100101100110,
64'b0000111111110000000011111111000001100110011001100110011001100110,
64'b0110100110010110011010011001011001011010101001011010010101011010,
64'b1111111100000000111111110000000010101010101010101010101010101010,
64'b1010101010101010101010101010101001100110011001100110011001100110,
64'b1001100101100110100110010110011001100110011001100110011001100110,
64'b0110100101101001100101101001011000001111000011111111000011110000,
64'b0000000011111111111111110000000001101001100101100110100110010110,
64'b1111000000001111000011111111000010101010101010101010101010101010,
64'b0000000011111111111111110000000011110000000011110000111111110000,
64'b1100110000110011001100111100110001101001011010011001011010010110,
64'b1010101001010101010101011010101011000011110000110011110000111100,
64'b1111000011110000111100001111000000000000111111111111111100000000,
64'b0110100110010110011010011001011011000011110000110011110000111100,
64'b1010101001010101010101011010101010010110100101101001011010010110,
64'b0011110011000011110000110011110011001100001100110011001111001100,
64'b0000000000000000000000000000000001100110011001100110011001100110,
64'b1100110011001100110011001100110010010110100101101001011010010110,
64'b1100001111000011001111000011110000111100001111000011110000111100,
64'b1100001100111100110000110011110011111111000000001111111100000000,
64'b0101010101010101101010101010101010010110011010010110100110010110,
64'b1010101001010101010101011010101011001100110011001100110011001100,
64'b0101010101010101101010101010101000000000111111111111111100000000,
64'b1010010110100101010110100101101001101001100101100110100110010110,
64'b1001100110011001011001100110011010100101010110101010010101011010,
64'b0101010110101010010101011010101001010101010101011010101010101010,
64'b0011110011000011110000110011110010100101010110101010010101011010,
64'b0011001100110011110011001100110001101001100101100110100110010110,
64'b0101101010100101101001010101101000001111000011111111000011110000,
64'b1010101010101010101010101010101010010110100101101001011010010110,
64'b0101101001011010010110100101101001101001100101100110100110010110,
64'b0000111111110000000011111111000000001111111100000000111111110000,
64'b0101101010100101101001010101101011111111111111110000000000000000,
64'b1100110011001100110011001100110000111100110000111100001100111100,
64'b1001100110011001011001100110011001011010010110100101101001011010,
64'b0110011001100110011001100110011011111111111111110000000000000000,
64'b1001100101100110100110010110011010010110011010010110100110010110,
64'b1001011010010110100101101001011011001100001100110011001111001100,
64'b1001100110011001011001100110011011001100110011001100110011001100,
64'b1111000000001111000011111111000001100110100110011001100101100110,
64'b0101101001011010010110100101101000111100110000111100001100111100,
64'b0110011010011001100110010110011011111111000000001111111100000000,
64'b0110011001100110011001100110011001101001100101100110100110010110,
64'b0101010101010101101010101010101001010101101010100101010110101010,
64'b0011110011000011110000110011110011000011001111001100001100111100,
64'b0000000000000000000000000000000010100101010110101010010101011010,
64'b0110011001100110011001100110011010010110100101101001011010010110,
64'b0011001111001100001100111100110011111111000000001111111100000000,
64'b0000111111110000000011111111000001011010101001011010010101011010,
64'b1010101001010101010101011010101011110000111100001111000011110000,
64'b0000000011111111111111110000000011111111111111110000000000000000,
64'b0011110011000011110000110011110011110000111100001111000011110000,
64'b0000000000000000000000000000000001100110011001100110011001100110,
64'b1111111111111111000000000000000011001100001100110011001111001100,
64'b0101010110101010010101011010101001101001100101100110100110010110,
64'b1010010101011010101001010101101000111100001111000011110000111100,
64'b0011001100110011110011001100110010011001100110010110011001100110,
64'b0110011001100110011001100110011011110000000011110000111111110000,
64'b1010101010101010101010101010101011001100001100110011001111001100,
64'b0101101001011010010110100101101011000011001111001100001100111100,
64'b0011110011000011110000110011110011111111111111110000000000000000,
64'b0000111100001111111100001111000011001100001100110011001111001100,
64'b1001100101100110100110010110011001010101101010100101010110101010,
64'b0101010110101010010101011010101000000000000000000000000000000000,
64'b0110011001100110011001100110011001010101101010100101010110101010,
64'b1010101010101010101010101010101000111100001111000011110000111100,
64'b1111111111111111000000000000000000001111000011111111000011110000,
64'b1100110000110011001100111100110010010110011010010110100110010110,
64'b1001011010010110100101101001011000001111111100000000111111110000,
64'b1010010110100101010110100101101000111100001111000011110000111100,
64'b1010101001010101010101011010101010101010010101010101010110101010,
64'b1100110011001100110011001100110010100101101001010101101001011010,
64'b0101010110101010010101011010101001011010101001011010010101011010,
64'b1100001111000011001111000011110000000000000000000000000000000000,
64'b0101101001011010010110100101101010100101101001010101101001011010,
64'b1100001100111100110000110011110010011001100110010110011001100110,
64'b0011001111001100001100111100110000000000000000000000000000000000,
64'b0000000011111111111111110000000000110011001100111100110011001100,
64'b1100110011001100110011001100110000001111111100000000111111110000,
64'b1111111111111111000000000000000011111111000000001111111100000000,
64'b1111000000001111000011111111000010010110011010010110100110010110,
64'b1100110011001100110011001100110001010101101010100101010110101010,
64'b1001100101100110100110010110011000001111111100000000111111110000,
64'b1001100110011001011001100110011000110011001100111100110011001100,
64'b0101101001011010010110100101101010011001011001101001100101100110,
64'b0011001100110011110011001100110001100110100110011001100101100110,
64'b0000111111110000000011111111000010101010101010101010101010101010,
64'b1001100101100110100110010110011000110011110011000011001111001100,
64'b1111000000001111000011111111000010010110100101101001011010010110,
64'b0000111100001111111100001111000010101010101010101010101010101010,
64'b1111111111111111000000000000000011110000111100001111000011110000,
64'b0101101001011010010110100101101010101010010101010101010110101010,
64'b0000000000000000000000000000000011111111111111110000000000000000,
64'b1010101001010101010101011010101000111100110000111100001100111100,
64'b0101101001011010010110100101101001100110011001100110011001100110,
64'b1001011010010110100101101001011010101010010101010101010110101010,
64'b0000000011111111111111110000000011110000111100001111000011110000,
64'b1001100101100110100110010110011001101001011010011001011010010110,
64'b1001011010010110100101101001011011000011110000110011110000111100,
64'b1001100110011001011001100110011001100110011001100110011001100110,
64'b1100110000110011001100111100110000001111000011111111000011110000,
64'b1010101010101010101010101010101011000011001111001100001100111100,
64'b0101010101010101101010101010101011001100110011001100110011001100,
64'b1001011001101001011010011001011011111111000000001111111100000000,
64'b1001100101100110100110010110011000110011001100111100110011001100,
64'b1111111111111111000000000000000010101010101010101010101010101010,
64'b0110011010011001100110010110011001011010101001011010010101011010,
64'b0011110000111100001111000011110010010110100101101001011010010110,
64'b0011110011000011110000110011110000110011001100111100110011001100,
64'b1100001100111100110000110011110001010101101010100101010110101010,
64'b0110100101101001100101101001011011000011001111001100001100111100,
64'b1010010101011010101001010101101010100101010110101010010101011010,
64'b0000111111110000000011111111000010010110100101101001011010010110,
64'b1010101001010101010101011010101011111111000000001111111100000000,
64'b1100110000110011001100111100110001011010101001011010010101011010,
64'b1100110000110011001100111100110011110000111100001111000011110000,
64'b1010101010101010101010101010101011111111111111110000000000000000,
64'b0110100101101001100101101001011011110000111100001111000011110000,
64'b1111111111111111000000000000000001100110011001100110011001100110,
64'b0011110011000011110000110011110011001100001100110011001111001100,
64'b0000000000000000000000000000000001101001100101100110100110010110,
64'b0101101010100101101001010101101010100101101001010101101001011010,
64'b0101101010100101101001010101101010100101010110101010010101011010,
64'b1100001100111100110000110011110011110000000011110000111111110000,
64'b0110011010011001100110010110011010101010010101010101010110101010,
64'b0000000011111111111111110000000011110000111100001111000011110000,
64'b0011001100110011110011001100110011110000000011110000111111110000,
64'b1010010110100101010110100101101001100110011001100110011001100110,
64'b1010010110100101010110100101101001010101010101011010101010101010,
64'b0110011001100110011001100110011000111100110000111100001100111100,
64'b1100001100111100110000110011110001010101101010100101010110101010,
64'b1010101010101010101010101010101011000011110000110011110000111100,
64'b0101101010100101101001010101101001011010101001011010010101011010,
64'b1010101010101010101010101010101011001100110011001100110011001100,
64'b0011001111001100001100111100110001100110100110011001100101100110,
64'b0101101001011010010110100101101001011010010110100101101001011010,
64'b0101101010100101101001010101101000000000111111111111111100000000,
64'b1010010110100101010110100101101011111111111111110000000000000000,
64'b0110011010011001100110010110011001100110011001100110011001100110,
64'b0101010110101010010101011010101000001111000011111111000011110000,
64'b0011001100110011110011001100110000111100110000111100001100111100,
64'b1001100110011001011001100110011011001100001100110011001111001100,
64'b1010101001010101010101011010101001100110011001100110011001100110,
64'b1111000000001111000011111111000010011001100110010110011001100110,
64'b0011001100110011110011001100110011110000000011110000111111110000,
64'b1001100110011001011001100110011000110011001100111100110011001100,
64'b1100001100111100110000110011110011111111000000001111111100000000,
64'b0101101001011010010110100101101001101001011010011001011010010110,
64'b0000111100001111111100001111000010011001011001101001100101100110,
64'b1100110000110011001100111100110011111111111111110000000000000000,
64'b1111111100000000111111110000000010101010101010101010101010101010,
64'b0101101010100101101001010101101010010110100101101001011010010110,
64'b1001011001101001011010011001011011111111000000001111111100000000,
64'b0101101010100101101001010101101001011010101001011010010101011010,
64'b1001011001101001011010011001011010100101101001010101101001011010,
64'b1010010101011010101001010101101010010110100101101001011010010110,
64'b1010101001010101010101011010101000111100001111000011110000111100,
64'b1010010110100101010110100101101010101010010101010101010110101010,
64'b1100001100111100110000110011110001011010010110100101101001011010,
64'b0000000000000000000000000000000010101010101010101010101010101010,
64'b0011001111001100001100111100110001101001100101100110100110010110,
64'b1111111100000000111111110000000001101001011010011001011010010110,
64'b1010010110100101010110100101101000000000000000000000000000000000,
64'b0101010101010101101010101010101001100110011001100110011001100110,
64'b1100110000110011001100111100110011000011001111001100001100111100,
64'b1001011001101001011010011001011011111111111111110000000000000000,
64'b0110011010011001100110010110011011001100001100110011001111001100,
64'b1001011001101001011010011001011010011001011001101001100101100110,
64'b0110011010011001100110010110011001101001100101100110100110010110,
64'b0011001100110011110011001100110000001111111100000000111111110000,
64'b1001100101100110100110010110011000110011001100111100110011001100,
64'b0101101010100101101001010101101010011001011001101001100101100110,
64'b0000000000000000000000000000000011001100110011001100110011001100,
64'b1111000011110000111100001111000001101001100101100110100110010110,
64'b1100001100111100110000110011110011111111111111110000000000000000,
64'b0011001111001100001100111100110010101010101010101010101010101010,
64'b0000000000000000000000000000000001011010010110100101101001011010,
64'b1001011001101001011010011001011011000011110000110011110000111100,
64'b1001100110011001011001100110011000001111111100000000111111110000,
64'b1100001100111100110000110011110000001111111100000000111111110000,
64'b1001011010010110100101101001011001101001100101100110100110010110,
64'b0101010110101010010101011010101000000000000000000000000000000000,
64'b0101101001011010010110100101101000000000111111111111111100000000,
64'b1001011010010110100101101001011000001111000011111111000011110000,
64'b1001100110011001011001100110011000111100110000111100001100111100,
64'b0000111111110000000011111111000001010101101010100101010110101010,
64'b0000000011111111111111110000000000111100110000111100001100111100,
64'b1100110011001100110011001100110000000000000000000000000000000000,
64'b0000111100001111111100001111000001100110011001100110011001100110,
64'b0110011001100110011001100110011000110011110011000011001111001100,
64'b0000111100001111111100001111000000001111111100000000111111110000,
64'b1001100101100110100110010110011010101010010101010101010110101010,
64'b1111000011110000111100001111000000000000111111111111111100000000,
64'b1100001111000011001111000011110000111100110000111100001100111100,
64'b0000111111110000000011111111000000000000000000000000000000000000,
64'b0011001111001100001100111100110011111111111111110000000000000000,
64'b0011110011000011110000110011110001010101101010100101010110101010,
64'b0110100110010110011010011001011001011010101001011010010101011010,
64'b1111000011110000111100001111000001100110011001100110011001100110,
64'b1010101010101010101010101010101001011010101001011010010101011010,
64'b0110011010011001100110010110011010101010101010101010101010101010,
64'b1111111100000000111111110000000000111100001111000011110000111100,
64'b1111000011110000111100001111000000001111000011111111000011110000,
64'b1100110011001100110011001100110000000000111111111111111100000000,
64'b0110011010011001100110010110011000110011001100111100110011001100,
64'b0101010101010101101010101010101001010101010101011010101010101010,
64'b0000111100001111111100001111000001011010101001011010010101011010,
64'b1001011010010110100101101001011010101010101010101010101010101010,
64'b0000111100001111111100001111000000000000000000000000000000000000,
64'b0000111111110000000011111111000010011001100110010110011001100110,
64'b1100001111000011001111000011110011001100001100110011001111001100,
64'b0101101001011010010110100101101010010110100101101001011010010110,
64'b0110011001100110011001100110011011001100001100110011001111001100,
64'b1100001111000011001111000011110001100110011001100110011001100110,
64'b0101010101010101101010101010101000001111111100000000111111110000,
64'b1111111100000000111111110000000011111111000000001111111100000000,
64'b1111000011110000111100001111000001010101010101011010101010101010,
64'b1100001111000011001111000011110001011010010110100101101001011010,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b0101010110101010010101011010101001100110100110011001100101100110,
64'b0110100110010110011010011001011001100110011001100110011001100110,
64'b1111111100000000111111110000000000000000000000000000000000000000,
64'b1010101001010101010101011010101000111100001111000011110000111100,
64'b0000111111110000000011111111000010100101101001010101101001011010,
64'b1001100101100110100110010110011001101001100101100110100110010110,
64'b0011110000111100001111000011110000001111000011111111000011110000,
64'b0000111111110000000011111111000010010110100101101001011010010110,
64'b0110011001100110011001100110011000000000111111111111111100000000,
64'b0101010101010101101010101010101011111111111111110000000000000000,
64'b1111111100000000111111110000000011001100110011001100110011001100,
64'b0000111111110000000011111111000010011001011001101001100101100110,
64'b1001011010010110100101101001011000111100001111000011110000111100,
64'b0011001100110011110011001100110011000011110000110011110000111100,
64'b0011110011000011110000110011110010010110100101101001011010010110,
64'b1111111111111111000000000000000000000000000000000000000000000000,
64'b0011001100110011110011001100110000001111111100000000111111110000,
64'b1010101001010101010101011010101000110011110011000011001111001100,
64'b0011110000111100001111000011110001101001100101100110100110010110,
64'b0000111111110000000011111111000011111111000000001111111100000000,
64'b0000000011111111111111110000000001101001100101100110100110010110,
64'b0011110000111100001111000011110011111111111111110000000000000000,
64'b1100110011001100110011001100110010101010101010101010101010101010,
64'b0101010101010101101010101010101001011010010110100101101001011010,
64'b0000000011111111111111110000000011000011110000110011110000111100,
64'b1100001100111100110000110011110000001111111100000000111111110000,
64'b1111000011110000111100001111000000001111111100000000111111110000,
64'b0101101010100101101001010101101001101001100101100110100110010110,
64'b1010101010101010101010101010101000000000000000000000000000000000,
64'b0101101001011010010110100101101000000000111111111111111100000000,
64'b1001100110011001011001100110011000001111000011111111000011110000,
64'b1010010101011010101001010101101011000011001111001100001100111100,
64'b1001011010010110100101101001011000110011001100111100110011001100,
64'b0110100101101001100101101001011000001111111100000000111111110000,
64'b0110011001100110011001100110011001010101101010100101010110101010,
64'b0110100110010110011010011001011010100101101001010101101001011010,
64'b1010010110100101010110100101101001010101010101011010101010101010,
64'b0000000000000000000000000000000000111100110000111100001100111100,
64'b0000111100001111111100001111000001100110011001100110011001100110,
64'b1001100101100110100110010110011001100110100110011001100101100110,
64'b1111000011110000111100001111000001100110011001100110011001100110,
64'b1010101010101010101010101010101010010110100101101001011010010110,
64'b1100110011001100110011001100110011001100001100110011001111001100,
64'b1100110011001100110011001100110010100101010110101010010101011010,
64'b0101010110101010010101011010101000000000000000000000000000000000,
64'b1111111100000000111111110000000011110000111100001111000011110000,
64'b1010101001010101010101011010101010101010010101010101010110101010,
64'b1111000011110000111100001111000000110011001100111100110011001100,
64'b0101010101010101101010101010101000110011110011000011001111001100,
64'b1001011001101001011010011001011001100110011001100110011001100110,
64'b1010101010101010101010101010101001011010101001011010010101011010,
64'b1111000000001111000011111111000010010110100101101001011010010110,
64'b1111000000001111000011111111000011000011110000110011110000111100,
64'b0000111111110000000011111111000010010110100101101001011010010110,
64'b0110011001100110011001100110011011000011001111001100001100111100,
64'b0011110000111100001111000011110000001111000011111111000011110000,
64'b0011110000111100001111000011110001100110100110011001100101100110,
64'b1001100101100110100110010110011000000000000000000000000000000000,
64'b0110100101101001100101101001011001010101101010100101010110101010,
64'b0101101001011010010110100101101000110011001100111100110011001100,
64'b0011001111001100001100111100110001011010010110100101101001011010,
64'b1010010101011010101001010101101010100101101001010101101001011010,
64'b0011001111001100001100111100110000111100001111000011110000111100,
64'b0110011001100110011001100110011011001100001100110011001111001100,
64'b0000111111110000000011111111000001101001100101100110100110010110,
64'b0011001100110011110011001100110000001111111100000000111111110000,
64'b0101101010100101101001010101101001101001100101100110100110010110,
64'b1001011010010110100101101001011011110000000011110000111111110000,
64'b1100001100111100110000110011110011111111000000001111111100000000,
64'b1100001100111100110000110011110001101001011010011001011010010110,
64'b0110100110010110011010011001011010101010101010101010101010101010,
64'b1100001100111100110000110011110010011001100110010110011001100110,
64'b1001100101100110100110010110011011110000111100001111000011110000,
64'b0000111100001111111100001111000010011001011001101001100101100110,
64'b1100110000110011001100111100110000110011110011000011001111001100,
64'b0000111100001111111100001111000010100101010110101010010101011010,
64'b0011110000111100001111000011110000001111000011111111000011110000,
64'b0000000011111111111111110000000010010110011010010110100110010110,
64'b1111000011110000111100001111000000000000111111111111111100000000,
64'b0110011010011001100110010110011000111100110000111100001100111100,
64'b0110100110010110011010011001011000000000111111111111111100000000,
64'b1111000000001111000011111111000001010101010101011010101010101010,
64'b1111000000001111000011111111000011000011001111001100001100111100,
64'b1100001100111100110000110011110001100110011001100110011001100110,
64'b0110011010011001100110010110011000111100001111000011110000111100,
64'b1010101010101010101010101010101001010101101010100101010110101010,
64'b1001100101100110100110010110011011000011110000110011110000111100,
64'b1100110000110011001100111100110000001111000011111111000011110000,
64'b1111000000001111000011111111000011001100001100110011001111001100,
64'b1010010101011010101001010101101011111111000000001111111100000000,
64'b1111000011110000111100001111000010010110011010010110100110010110,
64'b1100110011001100110011001100110001010101010101011010101010101010,
64'b0011001100110011110011001100110001011010101001011010010101011010,
64'b0011110011000011110000110011110001010101010101011010101010101010,
64'b1100110000110011001100111100110001100110011001100110011001100110,
64'b0110011010011001100110010110011001011010101001011010010101011010,
64'b1111000011110000111100001111000000111100001111000011110000111100,
64'b0101010101010101101010101010101000001111111100000000111111110000,
64'b0000111100001111111100001111000000110011001100111100110011001100,
64'b1010010110100101010110100101101000001111111100000000111111110000,
64'b0110011010011001100110010110011001010101101010100101010110101010,
64'b0000111111110000000011111111000010100101101001010101101001011010,
64'b0110011010011001100110010110011001010101010101011010101010101010,
64'b1111000000001111000011111111000000111100110000111100001100111100,
64'b0110100110010110011010011001011001100110011001100110011001100110,
64'b0000000000000000000000000000000001100110100110011001100101100110,
64'b1111000000001111000011111111000001100110011001100110011001100110,
64'b0110100101101001100101101001011010010110100101101001011010010110,
64'b1010010110100101010110100101101011001100001100110011001111001100,
64'b0000000000000000000000000000000010100101010110101010010101011010,
64'b1100110011001100110011001100110000111100110000111100001100111100,
64'b0101010110101010010101011010101010011001100110010110011001100110,
64'b1001100101100110100110010110011011001100001100110011001111001100,
64'b0110100101101001100101101001011001011010101001011010010101011010,
64'b1010101001010101010101011010101010010110011010010110100110010110,
64'b1100001111000011001111000011110001100110011001100110011001100110,
64'b1010101001010101010101011010101001010101101010100101010110101010,
64'b1001011001101001011010011001011000001111111100000000111111110000,
64'b0000000000000000000000000000000000110011001100111100110011001100,
64'b0000000011111111111111110000000000111100001111000011110000111100,
64'b0110100110010110011010011001011000001111111100000000111111110000,
64'b1001100101100110100110010110011011000011110000110011110000111100,
64'b1010101010101010101010101010101011001100110011001100110011001100,
64'b0110011001100110011001100110011001100110100110011001100101100110,
64'b0101101001011010010110100101101011111111111111110000000000000000,
64'b1010010110100101010110100101101011000011110000110011110000111100,
64'b1010101010101010101010101010101000001111000011111111000011110000,
64'b0011110000111100001111000011110000110011110011000011001111001100,
64'b1010010101011010101001010101101010010110100101101001011010010110,
64'b1001011010010110100101101001011000111100001111000011110000111100,
64'b0000111100001111111100001111000010011001100110010110011001100110,
64'b0101101001011010010110100101101000000000000000000000000000000000,
64'b0101010101010101101010101010101000001111111100000000111111110000,
64'b0101101010100101101001010101101011001100001100110011001111001100,
64'b0000111100001111111100001111000011000011001111001100001100111100,
64'b1001100101100110100110010110011000001111111100000000111111110000,
64'b0000000000000000000000000000000001101001011010011001011010010110,
64'b0101101010100101101001010101101010101010101010101010101010101010,
64'b0101010110101010010101011010101010100101010110101010010101011010,
64'b0000111111110000000011111111000001010101101010100101010110101010,
64'b1010101001010101010101011010101010100101101001010101101001011010,
64'b1100110000110011001100111100110011000011001111001100001100111100,
64'b1100110000110011001100111100110000001111111100000000111111110000,
64'b0110011001100110011001100110011000111100001111000011110000111100,
64'b0110100110010110011010011001011010101010101010101010101010101010,
64'b0110011001100110011001100110011000000000111111111111111100000000,
64'b1010101001010101010101011010101000001111000011111111000011110000,
64'b1001100101100110100110010110011001011010101001011010010101011010,
64'b1100001100111100110000110011110011111111000000001111111100000000,
64'b0000000000000000000000000000000011000011001111001100001100111100,
64'b1100110000110011001100111100110001100110011001100110011001100110,
64'b1001100110011001011001100110011011001100001100110011001111001100,
64'b0000000011111111111111110000000000110011001100111100110011001100,
64'b0011001100110011110011001100110000110011110011000011001111001100,
64'b1010010110100101010110100101101001011010101001011010010101011010,
64'b1010010110100101010110100101101000000000111111111111111100000000,
64'b1001011010010110100101101001011000001111111100000000111111110000,
64'b0011110011000011110000110011110011001100110011001100110011001100,
64'b0011110000111100001111000011110011111111111111110000000000000000,
64'b0011001100110011110011001100110001010101101010100101010110101010,
64'b0110100101101001100101101001011001100110100110011001100101100110,
64'b0000111111110000000011111111000010101010101010101010101010101010,
64'b1001011010010110100101101001011001100110100110011001100101100110,
64'b0110011001100110011001100110011001010101010101011010101010101010,
64'b1111000011110000111100001111000001101001011010011001011010010110,
64'b0011110011000011110000110011110000110011110011000011001111001100,
64'b1111111111111111000000000000000000000000000000000000000000000000,
64'b1001100101100110100110010110011011001100001100110011001111001100,
64'b1001011001101001011010011001011001011010010110100101101001011010,
64'b1111000011110000111100001111000000110011001100111100110011001100,
64'b0000000011111111111111110000000000000000000000000000000000000000,
64'b0000111111110000000011111111000010101010101010101010101010101010,
64'b0011110000111100001111000011110001010101010101011010101010101010,
64'b1010010101011010101001010101101000001111000011111111000011110000,
64'b0000000000000000000000000000000000110011110011000011001111001100,
64'b1111111100000000111111110000000001101001011010011001011010010110,
64'b0101010101010101101010101010101001100110011001100110011001100110,
64'b1001100101100110100110010110011001101001100101100110100110010110,
64'b1001100110011001011001100110011010100101101001010101101001011010,
64'b0000111100001111111100001111000000000000000000000000000000000000,
64'b0110100101101001100101101001011000001111000011111111000011110000,
64'b0011001111001100001100111100110010011001011001101001100101100110,
64'b1100110011001100110011001100110011110000111100001111000011110000,
64'b0000111100001111111100001111000010101010101010101010101010101010,
64'b0000000011111111111111110000000011001100110011001100110011001100,
64'b1100001100111100110000110011110011001100110011001100110011001100,
64'b0000000011111111111111110000000001010101101010100101010110101010,
64'b0101010110101010010101011010101001011010010110100101101001011010,
64'b0110100101101001100101101001011011000011001111001100001100111100,
64'b1010010110100101010110100101101010010110100101101001011010010110,
64'b0000111100001111111100001111000000111100110000111100001100111100,
64'b0101010110101010010101011010101000110011110011000011001111001100,
64'b1111000000001111000011111111000010101010101010101010101010101010,
64'b0110100110010110011010011001011011111111000000001111111100000000,
64'b1010101010101010101010101010101001101001011010011001011010010110,
64'b0110100110010110011010011001011011111111000000001111111100000000,
64'b0000111111110000000011111111000011001100110011001100110011001100,
64'b1111111111111111000000000000000011110000111100001111000011110000,
64'b1001011001101001011010011001011011110000111100001111000011110000,
64'b0011001100110011110011001100110000110011001100111100110011001100,
64'b0011001111001100001100111100110000110011110011000011001111001100,
64'b1100001100111100110000110011110011110000000011110000111111110000,
64'b1001100101100110100110010110011011000011001111001100001100111100,
64'b0101010110101010010101011010101011110000000011110000111111110000,
64'b1001100110011001011001100110011010100101101001010101101001011010,
64'b0000000011111111111111110000000011001100110011001100110011001100,
64'b1001011001101001011010011001011011111111111111110000000000000000,
64'b1100110011001100110011001100110011000011001111001100001100111100,
64'b0011110011000011110000110011110001010101010101011010101010101010,
64'b0000000011111111111111110000000011110000111100001111000011110000,
64'b0000000000000000000000000000000011111111000000001111111100000000,
64'b1001011001101001011010011001011011111111000000001111111100000000,
64'b0101101001011010010110100101101011110000111100001111000011110000,
64'b0101101001011010010110100101101001011010010110100101101001011010,
64'b0101101010100101101001010101101010101010010101010101010110101010,
64'b1100001111000011001111000011110001011010101001011010010101011010,
64'b0011001100110011110011001100110000000000111111111111111100000000,
64'b0011110000111100001111000011110010011001011001101001100101100110,
64'b0101010101010101101010101010101001011010010110100101101001011010,
64'b1001011001101001011010011001011000000000000000000000000000000000,
64'b0101101001011010010110100101101001011010101001011010010101011010,
64'b1111000000001111000011111111000011001100110011001100110011001100,
64'b0101010101010101101010101010101001010101101010100101010110101010,
64'b1010101010101010101010101010101011111111111111110000000000000000,
64'b0011110011000011110000110011110011111111111111110000000000000000,
64'b1001100101100110100110010110011011111111000000001111111100000000,
64'b0011001111001100001100111100110000110011110011000011001111001100,
64'b1100110000110011001100111100110010011001100110010110011001100110,
64'b1010010101011010101001010101101001100110100110011001100101100110,
64'b0101101001011010010110100101101001010101010101011010101010101010,
64'b1010010101011010101001010101101001101001011010011001011010010110,
64'b1100110011001100110011001100110000110011110011000011001111001100,
64'b1001011001101001011010011001011000000000000000000000000000000000,
64'b1001100101100110100110010110011011001100001100110011001111001100,
64'b0000000011111111111111110000000001011010010110100101101001011010,
64'b0110011001100110011001100110011000110011001100111100110011001100,
64'b0110011001100110011001100110011000000000000000000000000000000000,
64'b1111000000001111000011111111000010101010101010101010101010101010,
64'b0110100101101001100101101001011001010101010101011010101010101010,
64'b1111000011110000111100001111000011110000111100001111000011110000,
64'b0011001111001100001100111100110011111111111111110000000000000000,
64'b1010101001010101010101011010101000001111111100000000111111110000,
64'b0000111111110000000011111111000000001111000011111111000011110000,
64'b0000111111110000000011111111000011111111000000001111111100000000,
64'b1001100101100110100110010110011010101010101010101010101010101010,
64'b1111000011110000111100001111000010011001011001101001100101100110,
64'b0110100101101001100101101001011001101001011010011001011010010110,
64'b1100110000110011001100111100110011001100110011001100110011001100,
64'b1001011001101001011010011001011010010110011010010110100110010110,
64'b1100001111000011001111000011110001101001011010011001011010010110,
64'b0000000011111111111111110000000011001100110011001100110011001100,
64'b0011001100110011110011001100110000000000000000000000000000000000,
64'b1100001100111100110000110011110001010101101010100101010110101010,
64'b1001011001101001011010011001011000000000000000000000000000000000,
64'b1001100101100110100110010110011010101010010101010101010110101010,
64'b1010010110100101010110100101101011111111000000001111111100000000,
64'b0000111100001111111100001111000001010101010101011010101010101010,
64'b0101101010100101101001010101101011001100110011001100110011001100,
64'b0000111111110000000011111111000011000011110000110011110000111100,
64'b1010101001010101010101011010101011000011001111001100001100111100,
64'b0110100110010110011010011001011001011010010110100101101001011010,
64'b0000000000000000000000000000000000111100110000111100001100111100,
64'b0110011010011001100110010110011001101001100101100110100110010110,
64'b0101010110101010010101011010101001011010010110100101101001011010,
64'b0110100101101001100101101001011000000000000000000000000000000000,
64'b0110011001100110011001100110011011001100110011001100110011001100,
64'b1010010110100101010110100101101000000000000000000000000000000000,
64'b1100001100111100110000110011110000110011001100111100110011001100,
64'b0011110000111100001111000011110001010101010101011010101010101010,
64'b0101101001011010010110100101101011001100110011001100110011001100,
64'b1111111111111111000000000000000001011010010110100101101001011010,
64'b0101101010100101101001010101101000001111111100000000111111110000,
64'b0101101001011010010110100101101001011010101001011010010101011010,
64'b0101101001011010010110100101101000110011110011000011001111001100,
64'b1001011001101001011010011001011011110000000011110000111111110000,
64'b0000000000000000000000000000000010010110011010010110100110010110,
64'b1001100101100110100110010110011000110011110011000011001111001100,
64'b1111000000001111000011111111000000000000000000000000000000000000,
64'b0101010110101010010101011010101011110000111100001111000011110000,
64'b1001100101100110100110010110011000000000000000000000000000000000,
64'b0101101010100101101001010101101011110000111100001111000011110000,
64'b0000111111110000000011111111000001100110011001100110011001100110,
64'b0011001111001100001100111100110001011010010110100101101001011010,
64'b0000000000000000000000000000000000110011110011000011001111001100,
64'b0110011010011001100110010110011000000000111111111111111100000000,
64'b1001100101100110100110010110011011001100001100110011001111001100,
64'b0011001111001100001100111100110010100101101001010101101001011010,
64'b0011110011000011110000110011110000000000111111111111111100000000,
64'b1010101010101010101010101010101010010110011010010110100110010110,
64'b1100001111000011001111000011110010100101101001010101101001011010,
64'b0000000011111111111111110000000000000000000000000000000000000000,
64'b0110011001100110011001100110011011111111000000001111111100000000,
64'b0101101010100101101001010101101000000000000000000000000000000000,
64'b0110011001100110011001100110011011111111000000001111111100000000,
64'b1010010110100101010110100101101000111100001111000011110000111100,
64'b0000000011111111111111110000000000110011110011000011001111001100,
64'b1001100101100110100110010110011000001111000011111111000011110000,
64'b0011001100110011110011001100110011111111111111110000000000000000,
64'b0000000000000000000000000000000010100101101001010101101001011010,
64'b1100001100111100110000110011110010011001011001101001100101100110,
64'b0110011001100110011001100110011001010101010101011010101010101010,
64'b1010010110100101010110100101101010010110011010010110100110010110,
64'b0000111100001111111100001111000010011001011001101001100101100110,
64'b0110011001100110011001100110011010101010101010101010101010101010,
64'b0101010110101010010101011010101000000000000000000000000000000000,
64'b1111111111111111000000000000000000000000000000000000000000000000,
64'b0011110011000011110000110011110011111111111111110000000000000000,
64'b0011110000111100001111000011110000001111111100000000111111110000,
64'b0101101010100101101001010101101000001111000011111111000011110000,
64'b1111000000001111000011111111000011111111000000001111111100000000,
64'b0000000000000000000000000000000010101010101010101010101010101010,
64'b1100001111000011001111000011110010011001011001101001100101100110,
64'b0011110000111100001111000011110001101001011010011001011010010110,
64'b1010101001010101010101011010101011001100110011001100110011001100,
64'b1111000000001111000011111111000010010110011010010110100110010110,
64'b0101010101010101101010101010101001101001011010011001011010010110,
64'b1010010110100101010110100101101011001100110011001100110011001100,
64'b0000111111110000000011111111000000000000000000000000000000000000,
64'b0000000000000000000000000000000010011001011001101001100101100110,
64'b0101101010100101101001010101101010101010010101010101010110101010,
64'b1010010101011010101001010101101010100101101001010101101001011010,
64'b1100110000110011001100111100110011110000111100001111000011110000,
64'b1010101001010101010101011010101011001100001100110011001111001100,
64'b1010101010101010101010101010101000111100001111000011110000111100,
64'b0000111111110000000011111111000010101010101010101010101010101010,
64'b1010010101011010101001010101101000001111000011111111000011110000,
64'b0011001100110011110011001100110011001100001100110011001111001100,
64'b1010101001010101010101011010101011111111000000001111111100000000,
64'b0110011001100110011001100110011001101001011010011001011010010110,
64'b1001100101100110100110010110011001101001011010011001011010010110,
64'b0101010110101010010101011010101011000011001111001100001100111100,
64'b0011001111001100001100111100110011110000000011110000111111110000,
64'b0110011001100110011001100110011010011001011001101001100101100110,
64'b0110100101101001100101101001011010010110100101101001011010010110,
64'b0000000011111111111111110000000001011010010110100101101001011010,
64'b0000000011111111111111110000000010010110011010010110100110010110,
64'b1001011010010110100101101001011001010101101010100101010110101010,
64'b0110100110010110011010011001011010100101101001010101101001011010,
64'b0000000000000000000000000000000000110011001100111100110011001100,
64'b0110011010011001100110010110011000110011110011000011001111001100,
64'b0101101001011010010110100101101010010110100101101001011010010110,
64'b1001011001101001011010011001011011000011110000110011110000111100,
64'b1111000011110000111100001111000001011010101001011010010101011010,
64'b0000111111110000000011111111000001100110011001100110011001100110,
64'b1001011001101001011010011001011010101010010101010101010110101010,
64'b1001011001101001011010011001011001101001011010011001011010010110,
64'b1100110011001100110011001100110011000011001111001100001100111100,
64'b0101101010100101101001010101101000110011110011000011001111001100,
64'b1100110000110011001100111100110000111100110000111100001100111100,
64'b1001100101100110100110010110011010011001100110010110011001100110,
64'b0101010110101010010101011010101000110011110011000011001111001100,
64'b1100110000110011001100111100110001011010010110100101101001011010,
64'b0101010110101010010101011010101010100101101001010101101001011010,
64'b0101101010100101101001010101101011000011001111001100001100111100,
64'b0011110000111100001111000011110000001111111100000000111111110000,
64'b0110011010011001100110010110011001100110100110011001100101100110,
64'b0011110000111100001111000011110010010110100101101001011010010110,
64'b1001011001101001011010011001011010011001100110010110011001100110,
64'b1001011001101001011010011001011001101001100101100110100110010110,
64'b0101101001011010010110100101101001011010101001011010010101011010,
64'b1100110000110011001100111100110000001111000011111111000011110000,
64'b1010010110100101010110100101101011110000000011110000111111110000,
64'b0110100101101001100101101001011010010110100101101001011010010110,
64'b0011001100110011110011001100110010100101101001010101101001011010,
64'b0000111100001111111100001111000000110011110011000011001111001100,
64'b1001100110011001011001100110011000110011110011000011001111001100,
64'b1100110000110011001100111100110001011010101001011010010101011010,
64'b1010010101011010101001010101101000000000111111111111111100000000,
64'b1100001111000011001111000011110011000011110000110011110000111100,
64'b1010010101011010101001010101101001101001100101100110100110010110,
64'b1010010110100101010110100101101000001111111100000000111111110000,
64'b0011110000111100001111000011110000111100001111000011110000111100,
64'b1001011010010110100101101001011011000011110000110011110000111100,
64'b0000000011111111111111110000000001011010010110100101101001011010,
64'b0000000000000000000000000000000000110011001100111100110011001100,
64'b1001100101100110100110010110011010011001011001101001100101100110,
64'b0011001100110011110011001100110001011010101001011010010101011010,
64'b1001100110011001011001100110011001101001100101100110100110010110,
64'b0000000011111111111111110000000010011001011001101001100101100110,
64'b0110011001100110011001100110011000001111111100000000111111110000,
64'b0110011001100110011001100110011001010101101010100101010110101010,
64'b0011110011000011110000110011110010010110011010010110100110010110,
64'b0101101001011010010110100101101010101010101010101010101010101010,
64'b0000000000000000000000000000000010101010010101010101010110101010,
64'b0000111100001111111100001111000000001111111100000000111111110000,
64'b1100110011001100110011001100110000001111111100000000111111110000,
64'b1111000000001111000011111111000010011001011001101001100101100110,
64'b0011001111001100001100111100110011110000111100001111000011110000,
64'b0011001100110011110011001100110001101001011010011001011010010110,
64'b1001100110011001011001100110011011001100001100110011001111001100,
64'b0101101010100101101001010101101010010110011010010110100110010110,
64'b1100001100111100110000110011110011000011110000110011110000111100,
64'b0101010101010101101010101010101000000000111111111111111100000000,
64'b0011110011000011110000110011110000110011001100111100110011001100,
64'b1100001100111100110000110011110000111100110000111100001100111100,
64'b0101101001011010010110100101101001100110011001100110011001100110,
64'b1001100101100110100110010110011000110011001100111100110011001100,
64'b0101010101010101101010101010101010101010010101010101010110101010,
64'b0101010110101010010101011010101000000000111111111111111100000000,
64'b0000111100001111111100001111000011000011110000110011110000111100,
64'b0011110011000011110000110011110011111111000000001111111100000000,
64'b0000000000000000000000000000000011000011001111001100001100111100,
64'b1111111111111111000000000000000010100101101001010101101001011010,
64'b1010101010101010101010101010101010010110011010010110100110010110,
64'b1100110011001100110011001100110010100101010110101010010101011010,
64'b0000111100001111111100001111000001010101010101011010101010101010,
64'b0101101001011010010110100101101001011010010110100101101001011010,
64'b0110100110010110011010011001011001011010101001011010010101011010,
64'b1111000011110000111100001111000010010110100101101001011010010110,
64'b0110100101101001100101101001011001011010010110100101101001011010,
64'b1100110011001100110011001100110010011001100110010110011001100110,
64'b1001100110011001011001100110011001010101010101011010101010101010,
64'b1111111100000000111111110000000010100101010110101010010101011010,
64'b0101101010100101101001010101101001010101010101011010101010101010,
64'b1010101010101010101010101010101011110000000011110000111111110000,
64'b0000000000000000000000000000000000110011110011000011001111001100,
64'b0110011001100110011001100110011010010110011010010110100110010110,
64'b1111000011110000111100001111000001100110100110011001100101100110,
64'b1111111100000000111111110000000011001100110011001100110011001100,
64'b1001100101100110100110010110011010011001011001101001100101100110,
64'b0011110011000011110000110011110011001100001100110011001111001100,
64'b1111111100000000111111110000000001101001100101100110100110010110,
64'b1100001100111100110000110011110000110011110011000011001111001100,
64'b0101101001011010010110100101101000111100001111000011110000111100,
64'b0011110000111100001111000011110001100110011001100110011001100110,
64'b0101010101010101101010101010101001100110100110011001100101100110,
64'b1100110000110011001100111100110011001100110011001100110011001100,
64'b0110011001100110011001100110011010101010010101010101010110101010,
64'b0000000000000000000000000000000010100101101001010101101001011010,
64'b0011110000111100001111000011110000111100110000111100001100111100,
64'b1111111100000000111111110000000001101001011010011001011010010110,
64'b1111111111111111000000000000000001011010010110100101101001011010,
64'b1100001111000011001111000011110011000011110000110011110000111100,
64'b1111000000001111000011111111000000001111000011111111000011110000,
64'b1010101010101010101010101010101001101001100101100110100110010110,
64'b0101101010100101101001010101101010100101101001010101101001011010,
64'b0011001111001100001100111100110000001111111100000000111111110000,
64'b0000111111110000000011111111000000111100001111000011110000111100,
64'b1100110011001100110011001100110011000011110000110011110000111100,
64'b1010010110100101010110100101101001011010010110100101101001011010,
64'b1001011010010110100101101001011000110011001100111100110011001100,
64'b0000000000000000000000000000000010011001011001101001100101100110,
64'b0000111111110000000011111111000001011010101001011010010101011010,
64'b1111111111111111000000000000000001101001100101100110100110010110,
64'b0000000000000000000000000000000010011001011001101001100101100110,
64'b1010010101011010101001010101101000001111111100000000111111110000,
64'b1010101001010101010101011010101001010101101010100101010110101010,
64'b0110011001100110011001100110011001101001100101100110100110010110,
64'b1001011010010110100101101001011010011001100110010110011001100110,
64'b0000111111110000000011111111000000001111000011111111000011110000,
64'b0000000011111111111111110000000010101010101010101010101010101010,
64'b0101101010100101101001010101101001101001100101100110100110010110,
64'b1100001111000011001111000011110001101001100101100110100110010110,
64'b0101101010100101101001010101101011110000000011110000111111110000,
64'b1111111100000000111111110000000011111111000000001111111100000000,
64'b1111000000001111000011111111000001011010010110100101101001011010,
64'b0000111111110000000011111111000011001100001100110011001111001100,
64'b1100110000110011001100111100110000001111000011111111000011110000,
64'b0000111100001111111100001111000011001100110011001100110011001100,
64'b0011001111001100001100111100110000000000111111111111111100000000,
64'b1100110011001100110011001100110011000011001111001100001100111100,
64'b1111111100000000111111110000000010010110100101101001011010010110,
64'b0000111100001111111100001111000001010101101010100101010110101010,
64'b1111111100000000111111110000000001100110011001100110011001100110,
64'b0011110000111100001111000011110000111100110000111100001100111100,
64'b0110011010011001100110010110011000111100110000111100001100111100,
64'b0011110000111100001111000011110000000000111111111111111100000000,
64'b1010101001010101010101011010101001010101010101011010101010101010,
64'b1111000011110000111100001111000000110011110011000011001111001100,
64'b1010010110100101010110100101101000001111000011111111000011110000,
64'b1100001100111100110000110011110001010101101010100101010110101010,
64'b0101101010100101101001010101101001011010010110100101101001011010,
64'b1001011001101001011010011001011011111111111111110000000000000000,
64'b0011110000111100001111000011110010100101010110101010010101011010,
64'b0110100101101001100101101001011011000011001111001100001100111100,
64'b1111000011110000111100001111000000110011001100111100110011001100,
64'b0101010110101010010101011010101000111100001111000011110000111100,
64'b0101010101010101101010101010101011110000000011110000111111110000,
64'b0000000000000000000000000000000001011010101001011010010101011010,
64'b1111111111111111000000000000000001010101010101011010101010101010,
64'b1100110000110011001100111100110001100110011001100110011001100110,
64'b1010010110100101010110100101101010100101101001010101101001011010,
64'b0011110000111100001111000011110011111111000000001111111100000000,
64'b1001011010010110100101101001011010011001100110010110011001100110,
64'b1100001100111100110000110011110000110011110011000011001111001100,
64'b1010010110100101010110100101101000000000000000000000000000000000,
64'b0110100110010110011010011001011010011001011001101001100101100110,
64'b0110100110010110011010011001011011110000000011110000111111110000,
64'b0101010110101010010101011010101011110000111100001111000011110000,
64'b0011001100110011110011001100110010100101010110101010010101011010,
64'b1100110011001100110011001100110000000000111111111111111100000000,
64'b1010101010101010101010101010101001100110100110011001100101100110,
64'b0000000000000000000000000000000001100110011001100110011001100110,
64'b1010010110100101010110100101101010010110100101101001011010010110,
64'b1001100101100110100110010110011000110011110011000011001111001100,
64'b1010010101011010101001010101101001010101010101011010101010101010,
64'b1100001100111100110000110011110000111100001111000011110000111100,
64'b1111000000001111000011111111000010100101101001010101101001011010,
64'b0011001111001100001100111100110000000000000000000000000000000000,
64'b0110100110010110011010011001011000111100001111000011110000111100,
64'b1010101001010101010101011010101010101010010101010101010110101010,
64'b0011110011000011110000110011110001010101101010100101010110101010,
64'b1111000000001111000011111111000011001100001100110011001111001100,
64'b0000000011111111111111110000000011111111111111110000000000000000,
64'b0000111100001111111100001111000001101001011010011001011010010110,
64'b0101101010100101101001010101101010010110100101101001011010010110,
64'b1100110011001100110011001100110011000011001111001100001100111100,
64'b1001100101100110100110010110011000001111000011111111000011110000,
64'b1100001111000011001111000011110011001100110011001100110011001100,
64'b0011110000111100001111000011110010100101010110101010010101011010,
64'b0000111111110000000011111111000000110011110011000011001111001100,
64'b1001011001101001011010011001011010101010101010101010101010101010,
64'b0000111111110000000011111111000000001111111100000000111111110000,
64'b0000111100001111111100001111000000110011001100111100110011001100,
64'b0101010101010101101010101010101010011001100110010110011001100110,
64'b1010101010101010101010101010101000001111000011111111000011110000,
64'b0000111111110000000011111111000010101010101010101010101010101010,
64'b1001011001101001011010011001011001101001100101100110100110010110,
64'b0011110000111100001111000011110001101001100101100110100110010110,
64'b1010010101011010101001010101101011110000000011110000111111110000,
64'b0011001111001100001100111100110011111111000000001111111100000000,
64'b0000000000000000000000000000000001011010010110100101101001011010,
64'b0110100101101001100101101001011011001100001100110011001111001100,
64'b0000111111110000000011111111000000001111000011111111000011110000,
64'b0000111100001111111100001111000011001100110011001100110011001100,
64'b1001100101100110100110010110011011111111000000001111111100000000,
64'b0101010110101010010101011010101001100110011001100110011001100110,
64'b0110011001100110011001100110011010011001011001101001100101100110,
64'b0110011001100110011001100110011001010101010101011010101010101010,
64'b0000000011111111111111110000000000111100110000111100001100111100,
64'b0011110011000011110000110011110011111111000000001111111100000000,
64'b1010010101011010101001010101101001100110011001100110011001100110,
64'b1100110000110011001100111100110011111111111111110000000000000000,
64'b0000111100001111111100001111000010100101010110101010010101011010,
64'b0000000000000000000000000000000000111100001111000011110000111100,
64'b1100001100111100110000110011110011000011001111001100001100111100,
64'b1010101001010101010101011010101001011010101001011010010101011010,
64'b1111111100000000111111110000000001101001100101100110100110010110,
64'b1001011010010110100101101001011011001100110011001100110011001100,
64'b0000111100001111111100001111000000000000000000000000000000000000,
64'b0011001111001100001100111100110011001100001100110011001111001100,
64'b0011110011000011110000110011110011001100001100110011001111001100,
64'b1010010101011010101001010101101000000000000000000000000000000000,
64'b1001100101100110100110010110011010010110100101101001011010010110,
64'b0011110000111100001111000011110001100110100110011001100101100110,
64'b1111000000001111000011111111000011111111000000001111111100000000,
64'b1010010110100101010110100101101010010110100101101001011010010110,
64'b1010010101011010101001010101101000000000000000000000000000000000,
64'b0011110000111100001111000011110000111100001111000011110000111100,
64'b0011110000111100001111000011110011000011001111001100001100111100,
64'b0110011010011001100110010110011010100101101001010101101001011010,
64'b0000111111110000000011111111000000111100001111000011110000111100,
64'b1100001100111100110000110011110000000000000000000000000000000000,
64'b1010101001010101010101011010101000001111000011111111000011110000,
64'b1111000011110000111100001111000010100101101001010101101001011010,
64'b0011110000111100001111000011110010101010101010101010101010101010,
64'b0000000000000000000000000000000011000011001111001100001100111100,
64'b0101010101010101101010101010101011000011110000110011110000111100,
64'b1111111111111111000000000000000001010101010101011010101010101010,
64'b0110100101101001100101101001011011000011001111001100001100111100,
64'b0110100101101001100101101001011000000000000000000000000000000000,
64'b1100001111000011001111000011110000001111111100000000111111110000,
64'b0000000011111111111111110000000011110000000011110000111111110000,
64'b1111000000001111000011111111000000110011110011000011001111001100,
64'b1001100101100110100110010110011010100101010110101010010101011010,
64'b1111000000001111000011111111000000000000000000000000000000000000,
64'b0011001100110011110011001100110011111111000000001111111100000000,
64'b0101010110101010010101011010101010011001011001101001100101100110,
64'b0000111111110000000011111111000001100110011001100110011001100110,
64'b0000000000000000000000000000000011110000000011110000111111110000,
64'b1100110011001100110011001100110000001111111100000000111111110000,
64'b1010101010101010101010101010101001100110011001100110011001100110,
64'b0110100110010110011010011001011001011010101001011010010101011010,
64'b0110100110010110011010011001011000000000000000000000000000000000,
64'b1010010101011010101001010101101000000000111111111111111100000000,
64'b0101010101010101101010101010101000000000111111111111111100000000,
64'b1010101001010101010101011010101010100101101001010101101001011010,
64'b1001011010010110100101101001011000110011110011000011001111001100,
64'b0011110011000011110000110011110000111100001111000011110000111100,
64'b0101010110101010010101011010101011110000000011110000111111110000,
64'b1001100101100110100110010110011011000011001111001100001100111100,
64'b0101101001011010010110100101101001100110100110011001100101100110,
64'b1100001111000011001111000011110011000011001111001100001100111100,
64'b1010101001010101010101011010101011110000111100001111000011110000,
64'b0011001111001100001100111100110011000011001111001100001100111100,
64'b1100110011001100110011001100110000111100001111000011110000111100,
64'b0011001100110011110011001100110010100101010110101010010101011010,
64'b0000000000000000000000000000000000110011110011000011001111001100,
64'b1100001111000011001111000011110001011010010110100101101001011010,
64'b1010101001010101010101011010101010101010101010101010101010101010,
64'b1010010101011010101001010101101010010110100101101001011010010110,
64'b0110011010011001100110010110011000001111111100000000111111110000,
64'b1001011001101001011010011001011000000000111111111111111100000000,
64'b1100001100111100110000110011110001011010101001011010010101011010,
64'b0110100101101001100101101001011011000011110000110011110000111100,
64'b1100110000110011001100111100110001011010101001011010010101011010,
64'b1100001100111100110000110011110011111111000000001111111100000000,
64'b0101101010100101101001010101101011110000000011110000111111110000,
64'b0000000011111111111111110000000000001111111100000000111111110000,
64'b1111111100000000111111110000000011001100001100110011001111001100,
64'b0110011010011001100110010110011000001111000011111111000011110000,
64'b0000000011111111111111110000000000110011110011000011001111001100,
64'b1010101001010101010101011010101011001100110011001100110011001100,
64'b0101010110101010010101011010101011000011001111001100001100111100,
64'b0101010101010101101010101010101000000000111111111111111100000000,
64'b1001100110011001011001100110011011111111111111110000000000000000,
64'b0101101001011010010110100101101001100110100110011001100101100110,
64'b1001100110011001011001100110011010100101010110101010010101011010,
64'b0110011001100110011001100110011001100110100110011001100101100110,
64'b0000000000000000000000000000000001010101010101011010101010101010,
64'b0011001100110011110011001100110000000000111111111111111100000000,
64'b1010010101011010101001010101101010101010010101010101010110101010,
64'b0101101010100101101001010101101000001111000011111111000011110000,
64'b0000111111110000000011111111000001010101101010100101010110101010,
64'b0101101001011010010110100101101010100101101001010101101001011010,
64'b1010101001010101010101011010101011110000111100001111000011110000,
64'b1010101010101010101010101010101000001111111100000000111111110000,
64'b1100110011001100110011001100110011111111111111110000000000000000,
64'b1001011010010110100101101001011010101010101010101010101010101010,
64'b1001100101100110100110010110011001101001011010011001011010010110,
64'b0011110000111100001111000011110001100110100110011001100101100110,
64'b1001011010010110100101101001011011000011110000110011110000111100,
64'b0000000000000000000000000000000001100110011001100110011001100110,
64'b1111000011110000111100001111000001010101010101011010101010101010,
64'b0110011010011001100110010110011010011001100110010110011001100110,
64'b1100110000110011001100111100110001010101101010100101010110101010,
64'b1010101001010101010101011010101010011001100110010110011001100110,
64'b0011001111001100001100111100110000110011110011000011001111001100,
64'b0011001100110011110011001100110001010101101010100101010110101010,
64'b0110011001100110011001100110011011111111000000001111111100000000,
64'b0101101001011010010110100101101010101010101010101010101010101010,
64'b1100001100111100110000110011110001100110011001100110011001100110,
64'b1100001111000011001111000011110011000011001111001100001100111100,
64'b0000111111110000000011111111000001101001011010011001011010010110,
64'b1100001100111100110000110011110010100101010110101010010101011010,
64'b0000000000000000000000000000000010010110100101101001011010010110,
64'b1111111100000000111111110000000011001100110011001100110011001100,
64'b1100001111000011001111000011110010010110100101101001011010010110,
64'b1010010110100101010110100101101010011001100110010110011001100110,
64'b1001100110011001011001100110011000111100001111000011110000111100,
64'b1010010110100101010110100101101010100101101001010101101001011010,
64'b1111000011110000111100001111000000110011001100111100110011001100,
64'b1001011010010110100101101001011000000000000000000000000000000000,
64'b0011001111001100001100111100110001100110011001100110011001100110,
64'b1111000000001111000011111111000000111100001111000011110000111100,
64'b0000111111110000000011111111000011110000000011110000111111110000,
64'b1010101001010101010101011010101011000011001111001100001100111100,
64'b1111000000001111000011111111000001100110100110011001100101100110,
64'b0000000000000000000000000000000011000011001111001100001100111100,
64'b1111111111111111000000000000000011110000111100001111000011110000,
64'b0000111111110000000011111111000011000011001111001100001100111100,
64'b1001100101100110100110010110011000111100001111000011110000111100,
64'b1001011010010110100101101001011010100101010110101010010101011010,
64'b1001100101100110100110010110011000110011110011000011001111001100,
64'b0101010110101010010101011010101001011010010110100101101001011010,
64'b1100001100111100110000110011110010101010101010101010101010101010,
64'b1111000000001111000011111111000010100101010110101010010101011010,
64'b0011110011000011110000110011110010101010010101010101010110101010,
64'b0000111100001111111100001111000000111100001111000011110000111100,
64'b0110011001100110011001100110011000000000000000000000000000000000,
64'b0110011010011001100110010110011010010110011010010110100110010110,
64'b0101010110101010010101011010101000111100110000111100001100111100,
64'b1010010110100101010110100101101010010110100101101001011010010110,
64'b0101010110101010010101011010101011000011110000110011110000111100,
64'b1010101010101010101010101010101001010101101010100101010110101010,
64'b1111111111111111000000000000000001011010101001011010010101011010,
64'b1010010101011010101001010101101000001111111100000000111111110000,
64'b0000000000000000000000000000000010010110100101101001011010010110,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b1111000011110000111100001111000001100110100110011001100101100110,
64'b0110011001100110011001100110011000110011001100111100110011001100,
64'b0101101010100101101001010101101010100101010110101010010101011010,
64'b1111000011110000111100001111000000000000000000000000000000000000,
64'b1010010101011010101001010101101000111100110000111100001100111100,
64'b1100110000110011001100111100110001011010101001011010010101011010,
64'b1001011001101001011010011001011001101001100101100110100110010110,
64'b1100110000110011001100111100110000001111111100000000111111110000,
64'b0110011001100110011001100110011010011001100110010110011001100110,
64'b1111111111111111000000000000000011001100001100110011001111001100,
64'b1100001111000011001111000011110010101010010101010101010110101010,
64'b0000000000000000000000000000000011000011001111001100001100111100,
64'b0110011001100110011001100110011011001100110011001100110011001100,
64'b0000111100001111111100001111000001101001011010011001011010010110,
64'b0000000011111111111111110000000001011010010110100101101001011010,
64'b1100001100111100110000110011110001100110100110011001100101100110,
64'b0011001111001100001100111100110000000000000000000000000000000000,
64'b1010101010101010101010101010101011110000000011110000111111110000,
64'b0101101010100101101001010101101001100110100110011001100101100110,
64'b0011001111001100001100111100110010010110011010010110100110010110,
64'b1111000000001111000011111111000000000000111111111111111100000000,
64'b0011110000111100001111000011110000111100001111000011110000111100,
64'b1111111111111111000000000000000010100101101001010101101001011010,
64'b0000000000000000000000000000000010011001100110010110011001100110,
64'b1010101010101010101010101010101001011010101001011010010101011010,
64'b1001011010010110100101101001011011110000111100001111000011110000,
64'b0101010110101010010101011010101001101001100101100110100110010110,
64'b0101010101010101101010101010101010011001011001101001100101100110,
64'b0101101010100101101001010101101011000011110000110011110000111100,
64'b0000111100001111111100001111000010101010101010101010101010101010,
64'b1100110011001100110011001100110000000000111111111111111100000000,
64'b1100110000110011001100111100110001101001011010011001011010010110,
64'b1010010110100101010110100101101010010110011010010110100110010110,
64'b0000000011111111111111110000000001010101010101011010101010101010,
64'b1010010101011010101001010101101010100101010110101010010101011010,
64'b0000000000000000000000000000000000110011110011000011001111001100,
64'b1010101010101010101010101010101010010110100101101001011010010110,
64'b1100110011001100110011001100110001100110100110011001100101100110,
64'b1100001100111100110000110011110001010101101010100101010110101010,
64'b0110100110010110011010011001011000111100110000111100001100111100,
64'b1111000000001111000011111111000011000011110000110011110000111100,
64'b0110100110010110011010011001011000001111111100000000111111110000,
64'b0011001111001100001100111100110001100110011001100110011001100110,
64'b0011110011000011110000110011110011111111111111110000000000000000,
64'b0101101010100101101001010101101001101001100101100110100110010110,
64'b0011110011000011110000110011110010010110011010010110100110010110,
64'b0000000011111111111111110000000001100110011001100110011001100110,
64'b1100110000110011001100111100110001100110100110011001100101100110,
64'b1111111111111111000000000000000000001111000011111111000011110000,
64'b0110100110010110011010011001011011000011001111001100001100111100,
64'b1111000011110000111100001111000011000011110000110011110000111100,
64'b1010010101011010101001010101101001100110011001100110011001100110,
64'b0110011001100110011001100110011001011010101001011010010101011010,
64'b0011110000111100001111000011110010100101010110101010010101011010,
64'b1001100101100110100110010110011010101010010101010101010110101010,
64'b0110100101101001100101101001011000111100001111000011110000111100,
64'b1001011010010110100101101001011000000000000000000000000000000000,
64'b0011001100110011110011001100110010010110011010010110100110010110,
64'b1111111100000000111111110000000000111100110000111100001100111100,
64'b0000000011111111111111110000000010010110100101101001011010010110,
64'b0000111100001111111100001111000011000011110000110011110000111100,
64'b0101010101010101101010101010101001010101101010100101010110101010,
64'b0011001100110011110011001100110001011010101001011010010101011010,
64'b1111111100000000111111110000000000001111111100000000111111110000,
64'b1001100101100110100110010110011010010110100101101001011010010110,
64'b1001011010010110100101101001011010010110100101101001011010010110,
64'b0000111111110000000011111111000001011010010110100101101001011010,
64'b1100001111000011001111000011110000111100001111000011110000111100,
64'b1100001100111100110000110011110011000011001111001100001100111100,
64'b0110100110010110011010011001011001100110100110011001100101100110,
64'b1111000011110000111100001111000001101001011010011001011010010110,
64'b0101010101010101101010101010101011111111000000001111111100000000,
64'b1111111111111111000000000000000000111100001111000011110000111100,
64'b0101010110101010010101011010101010100101010110101010010101011010,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b0101101001011010010110100101101001101001011010011001011010010110,
64'b0101010101010101101010101010101010101010010101010101010110101010,
64'b0011110000111100001111000011110001101001100101100110100110010110,
64'b0011001100110011110011001100110000110011001100111100110011001100,
64'b0011110000111100001111000011110000001111000011111111000011110000,
64'b0000000011111111111111110000000000000000111111111111111100000000,
64'b0011110011000011110000110011110010010110011010010110100110010110,
64'b0101101001011010010110100101101010100101010110101010010101011010,
64'b1010101010101010101010101010101000111100001111000011110000111100,
64'b0110100101101001100101101001011011110000111100001111000011110000,
64'b1111111100000000111111110000000001011010010110100101101001011010,
64'b0011001100110011110011001100110001100110100110011001100101100110,
64'b1100001111000011001111000011110011000011110000110011110000111100,
64'b1001011010010110100101101001011001100110011001100110011001100110,
64'b1100110011001100110011001100110010011001100110010110011001100110,
64'b0000111111110000000011111111000011000011001111001100001100111100,
64'b1010101001010101010101011010101011110000111100001111000011110000,
64'b1001100110011001011001100110011001010101101010100101010110101010,
64'b1111000011110000111100001111000001010101010101011010101010101010,
64'b0011110011000011110000110011110010010110011010010110100110010110,
64'b1111111111111111000000000000000001100110100110011001100101100110,
64'b1001100101100110100110010110011000001111111100000000111111110000,
64'b0110011010011001100110010110011011111111000000001111111100000000,
64'b0000000011111111111111110000000000110011110011000011001111001100,
64'b0101101001011010010110100101101011000011110000110011110000111100,
64'b0101101010100101101001010101101010100101010110101010010101011010,
64'b1100110011001100110011001100110010010110100101101001011010010110,
64'b1111000011110000111100001111000000111100001111000011110000111100,
64'b0101010110101010010101011010101010100101010110101010010101011010,
64'b1001100110011001011001100110011001010101101010100101010110101010,
64'b1001011010010110100101101001011000110011001100111100110011001100,
64'b0101010110101010010101011010101011001100110011001100110011001100,
64'b1111000000001111000011111111000010010110011010010110100110010110,
64'b1010101010101010101010101010101001101001011010011001011010010110,
64'b0110100101101001100101101001011010101010010101010101010110101010,
64'b1100001111000011001111000011110011111111111111110000000000000000,
64'b0101010101010101101010101010101000001111000011111111000011110000,
64'b1001100101100110100110010110011000001111111100000000111111110000,
64'b1100110000110011001100111100110001100110100110011001100101100110,
64'b0101101001011010010110100101101011000011001111001100001100111100,
64'b1111111100000000111111110000000000001111111100000000111111110000,
64'b1100110011001100110011001100110000110011110011000011001111001100,
64'b1100110000110011001100111100110001101001100101100110100110010110,
64'b0101010101010101101010101010101011001100001100110011001111001100,
64'b0011110000111100001111000011110001010101010101011010101010101010,
64'b0110011010011001100110010110011001011010101001011010010101011010,
64'b0000000011111111111111110000000000001111000011111111000011110000,
64'b1001011010010110100101101001011011001100001100110011001111001100,
64'b0000000011111111111111110000000000001111000011111111000011110000,
64'b0011001111001100001100111100110000000000000000000000000000000000,
64'b1100001111000011001111000011110000000000111111111111111100000000,
64'b1111000011110000111100001111000000111100001111000011110000111100,
64'b0011110000111100001111000011110011111111111111110000000000000000,
64'b1111111111111111000000000000000000000000111111111111111100000000,
64'b0101101001011010010110100101101001011010010110100101101001011010,
64'b0101010110101010010101011010101000111100110000111100001100111100,
64'b0101101010100101101001010101101000001111000011111111000011110000,
64'b1010101001010101010101011010101001100110011001100110011001100110,
64'b1010010110100101010110100101101001100110100110011001100101100110,
64'b0011001111001100001100111100110001010101101010100101010110101010,
64'b0011110000111100001111000011110010100101101001010101101001011010,
64'b0101101001011010010110100101101001010101101010100101010110101010,
64'b1111000000001111000011111111000010101010101010101010101010101010,
64'b1010010101011010101001010101101011111111111111110000000000000000,
64'b1010101001010101010101011010101010100101010110101010010101011010,
64'b1010101010101010101010101010101000000000000000000000000000000000,
64'b0000000000000000000000000000000001010101010101011010101010101010,
64'b0011001111001100001100111100110010011001011001101001100101100110,
64'b0110100110010110011010011001011001011010101001011010010101011010,
64'b1111000011110000111100001111000001010101101010100101010110101010,
64'b1001011010010110100101101001011010010110100101101001011010010110,
64'b1111111100000000111111110000000011000011110000110011110000111100,
64'b1100001100111100110000110011110010011001100110010110011001100110,
64'b0101101001011010010110100101101000110011110011000011001111001100,
64'b1001011001101001011010011001011010011001100110010110011001100110,
64'b0101010101010101101010101010101011001100110011001100110011001100,
64'b1100110000110011001100111100110000000000000000000000000000000000,
64'b1100110011001100110011001100110001100110100110011001100101100110,
64'b1100001100111100110000110011110000000000000000000000000000000000,
64'b0000000000000000000000000000000011001100110011001100110011001100,
64'b0101101001011010010110100101101010010110100101101001011010010110,
64'b0011110011000011110000110011110001100110100110011001100101100110,
64'b1111111100000000111111110000000010011001100110010110011001100110,
64'b1100001100111100110000110011110011000011001111001100001100111100,
64'b1111111111111111000000000000000000001111111100000000111111110000,
64'b1111000000001111000011111111000010010110100101101001011010010110,
64'b0011001111001100001100111100110010100101101001010101101001011010,
64'b0011110011000011110000110011110000111100001111000011110000111100,
64'b0110011001100110011001100110011001011010010110100101101001011010,
64'b1010010110100101010110100101101000000000000000000000000000000000,
64'b0101101001011010010110100101101011000011110000110011110000111100,
64'b1111000000001111000011111111000010101010101010101010101010101010,
64'b0000000000000000000000000000000011110000111100001111000011110000,
64'b0011001111001100001100111100110011000011001111001100001100111100,
64'b1111000000001111000011111111000001101001011010011001011010010110,
64'b0101010101010101101010101010101010010110100101101001011010010110,
64'b1111000000001111000011111111000001011010101001011010010101011010,
64'b0000000000000000000000000000000000000000111111111111111100000000,
64'b1010101001010101010101011010101011000011001111001100001100111100,
64'b1010010110100101010110100101101000110011110011000011001111001100,
64'b1111000000001111000011111111000010100101010110101010010101011010,
64'b1001011010010110100101101001011000110011110011000011001111001100,
64'b0011001111001100001100111100110000000000000000000000000000000000,
64'b1001100101100110100110010110011000001111111100000000111111110000,
64'b0000000011111111111111110000000001100110011001100110011001100110,
64'b1010101010101010101010101010101011111111000000001111111100000000,
64'b1111000011110000111100001111000000001111111100000000111111110000,
64'b0000000011111111111111110000000011000011001111001100001100111100,
64'b0110011001100110011001100110011001101001100101100110100110010110,
64'b1010101001010101010101011010101011001100001100110011001111001100,
64'b1010101010101010101010101010101001010101010101011010101010101010,
64'b0011001100110011110011001100110001011010101001011010010101011010,
64'b1001100101100110100110010110011000001111000011111111000011110000,
64'b1010101001010101010101011010101011001100001100110011001111001100,
64'b0110100110010110011010011001011000001111000011111111000011110000,
64'b0000111100001111111100001111000000000000000000000000000000000000,
64'b1100001111000011001111000011110000000000111111111111111100000000,
64'b1111111111111111000000000000000000111100001111000011110000111100,
64'b0110011001100110011001100110011011111111111111110000000000000000,
64'b1111111100000000111111110000000011111111000000001111111100000000,
64'b0110100101101001100101101001011000110011001100111100110011001100,
64'b0000000000000000000000000000000011000011110000110011110000111100,
64'b1010101001010101010101011010101001100110011001100110011001100110,
64'b0011110000111100001111000011110011111111000000001111111100000000,
64'b1010010110100101010110100101101011111111111111110000000000000000,
64'b0000000011111111111111110000000000111100001111000011110000111100,
64'b0011110011000011110000110011110000110011001100111100110011001100,
64'b0101010110101010010101011010101001010101101010100101010110101010,
64'b1001011001101001011010011001011011001100110011001100110011001100,
64'b1001011010010110100101101001011010010110011010010110100110010110,
64'b1111000000001111000011111111000011001100001100110011001111001100,
64'b0000000011111111111111110000000000111100110000111100001100111100,
64'b1010010101011010101001010101101011001100110011001100110011001100,
64'b1010101001010101010101011010101011110000111100001111000011110000,
64'b1010101010101010101010101010101010100101010110101010010101011010,
64'b1001100101100110100110010110011010010110100101101001011010010110,
64'b1001100101100110100110010110011011111111111111110000000000000000,
64'b1001011001101001011010011001011000000000000000000000000000000000,
64'b0101010110101010010101011010101010100101010110101010010101011010,
64'b0110011001100110011001100110011011110000111100001111000011110000,
64'b1100110000110011001100111100110010011001100110010110011001100110,
64'b1010101010101010101010101010101011110000111100001111000011110000,
64'b1111111100000000111111110000000000111100110000111100001100111100,
64'b1111000011110000111100001111000010100101101001010101101001011010,
64'b0101010110101010010101011010101001011010101001011010010101011010,
64'b0011110000111100001111000011110001011010010110100101101001011010,
64'b0101101001011010010110100101101011111111000000001111111100000000,
64'b0110011001100110011001100110011011001100001100110011001111001100,
64'b0110100110010110011010011001011011000011001111001100001100111100,
64'b1111111111111111000000000000000000000000000000000000000000000000,
64'b1001100101100110100110010110011010101010101010101010101010101010,
64'b1001100101100110100110010110011011001100001100110011001111001100,
64'b0000000011111111111111110000000011111111000000001111111100000000,
64'b0101101010100101101001010101101000111100001111000011110000111100,
64'b1111000000001111000011111111000001010101101010100101010110101010,
64'b0110100101101001100101101001011011110000000011110000111111110000,
64'b0000111100001111111100001111000010011001011001101001100101100110,
64'b0011001111001100001100111100110001100110100110011001100101100110,
64'b1010101010101010101010101010101010011001011001101001100101100110,
64'b0011001111001100001100111100110011111111111111110000000000000000,
64'b0011110000111100001111000011110000001111000011111111000011110000,
64'b0011110011000011110000110011110001011010101001011010010101011010,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0110100101101001100101101001011011001100110011001100110011001100,
64'b1100001111000011001111000011110000001111000011111111000011110000,
64'b1111111111111111000000000000000001010101010101011010101010101010,
64'b0110011010011001100110010110011000001111111100000000111111110000,
64'b1010101001010101010101011010101000110011001100111100110011001100,
64'b0110100110010110011010011001011000000000111111111111111100000000,
64'b0101010110101010010101011010101001101001011010011001011010010110,
64'b1010010110100101010110100101101011000011110000110011110000111100,
64'b1100110011001100110011001100110010010110100101101001011010010110,
64'b1100110011001100110011001100110010101010101010101010101010101010,
64'b0000111111110000000011111111000001010101101010100101010110101010,
64'b0101101001011010010110100101101001100110100110011001100101100110,
64'b1001011010010110100101101001011010101010101010101010101010101010,
64'b0110011010011001100110010110011011110000111100001111000011110000,
64'b1010010110100101010110100101101011111111000000001111111100000000,
64'b1001011001101001011010011001011001100110011001100110011001100110,
64'b0011110011000011110000110011110010101010010101010101010110101010,
64'b0000111111110000000011111111000011110000111100001111000011110000,
64'b0000000011111111111111110000000001010101010101011010101010101010,
64'b1100001100111100110000110011110001101001100101100110100110010110,
64'b0011001100110011110011001100110010100101010110101010010101011010,
64'b1111111100000000111111110000000001101001100101100110100110010110,
64'b0011001100110011110011001100110011001100110011001100110011001100,
64'b0000000011111111111111110000000000110011001100111100110011001100,
64'b1001100110011001011001100110011011000011110000110011110000111100,
64'b1111111100000000111111110000000001100110011001100110011001100110,
64'b0110011001100110011001100110011011111111000000001111111100000000,
64'b1001100110011001011001100110011011111111111111110000000000000000,
64'b1010101010101010101010101010101000111100001111000011110000111100,
64'b0000111100001111111100001111000000110011001100111100110011001100,
64'b0011110000111100001111000011110001010101101010100101010110101010,
64'b0110100101101001100101101001011011001100110011001100110011001100,
64'b1010101010101010101010101010101010010110011010010110100110010110,
64'b1111000000001111000011111111000011001100001100110011001111001100,
64'b0000111111110000000011111111000011000011001111001100001100111100,
64'b0101101001011010010110100101101010011001100110010110011001100110,
64'b0101010101010101101010101010101011110000111100001111000011110000,
64'b1001011010010110100101101001011000001111000011111111000011110000,
64'b0101010101010101101010101010101010101010101010101010101010101010,
64'b0011110000111100001111000011110001011010010110100101101001011010,
64'b0011110000111100001111000011110000000000111111111111111100000000,
64'b0110011001100110011001100110011010011001100110010110011001100110,
64'b1111111100000000111111110000000010100101010110101010010101011010,
64'b1010010101011010101001010101101000001111111100000000111111110000,
64'b1100001100111100110000110011110001100110011001100110011001100110,
64'b0110011001100110011001100110011011001100110011001100110011001100,
64'b0000000011111111111111110000000010100101010110101010010101011010,
64'b0101010110101010010101011010101000000000000000000000000000000000,
64'b0101101010100101101001010101101011111111111111110000000000000000,
64'b1100110011001100110011001100110001010101101010100101010110101010,
64'b1100001111000011001111000011110001010101010101011010101010101010,
64'b1111000011110000111100001111000001011010010110100101101001011010,
64'b0000000011111111111111110000000010010110011010010110100110010110,
64'b0000111100001111111100001111000011111111000000001111111100000000,
64'b0000000011111111111111110000000010101010010101010101010110101010,
64'b1010101001010101010101011010101000110011001100111100110011001100,
64'b0101101001011010010110100101101010010110100101101001011010010110,
64'b0110011010011001100110010110011010101010101010101010101010101010,
64'b1100110000110011001100111100110000000000111111111111111100000000,
64'b1111111100000000111111110000000011001100110011001100110011001100,
64'b1100001100111100110000110011110010100101010110101010010101011010,
64'b0000111111110000000011111111000010101010101010101010101010101010,
64'b0101101001011010010110100101101010011001100110010110011001100110,
64'b1010010110100101010110100101101011001100110011001100110011001100,
64'b0110100110010110011010011001011010011001011001101001100101100110,
64'b0101101001011010010110100101101000111100110000111100001100111100,
64'b0101010101010101101010101010101001010101010101011010101010101010,
64'b0110100110010110011010011001011000110011001100111100110011001100,
64'b1100110000110011001100111100110001011010010110100101101001011010,
64'b0000111100001111111100001111000001101001100101100110100110010110,
64'b0101010101010101101010101010101011001100110011001100110011001100,
64'b0101010110101010010101011010101011111111111111110000000000000000,
64'b0101010110101010010101011010101001011010010110100101101001011010,
64'b1010101010101010101010101010101000110011110011000011001111001100,
64'b1010101001010101010101011010101001100110011001100110011001100110,
64'b0011001111001100001100111100110000111100001111000011110000111100,
64'b0011001111001100001100111100110001011010010110100101101001011010,
64'b1001011001101001011010011001011011000011110000110011110000111100,
64'b0011001111001100001100111100110011110000000011110000111111110000,
64'b1100110011001100110011001100110001100110011001100110011001100110,
64'b1001011001101001011010011001011001011010010110100101101001011010,
64'b0000111100001111111100001111000010011001011001101001100101100110,
64'b0101010110101010010101011010101000111100110000111100001100111100,
64'b0110011001100110011001100110011011110000111100001111000011110000,
64'b1001100110011001011001100110011000000000000000000000000000000000,
64'b0011001100110011110011001100110010011001011001101001100101100110,
64'b1100110011001100110011001100110011110000111100001111000011110000,
64'b0101101001011010010110100101101011111111111111110000000000000000,
64'b1010010110100101010110100101101000001111111100000000111111110000,
64'b1010010101011010101001010101101010011001100110010110011001100110,
64'b0000000011111111111111110000000000110011110011000011001111001100,
64'b0000000000000000000000000000000000001111111100000000111111110000,
64'b1111000000001111000011111111000010010110011010010110100110010110,
64'b0000000000000000000000000000000000001111000011111111000011110000,
64'b0000000000000000000000000000000010010110011010010110100110010110,
64'b0000111111110000000011111111000001100110011001100110011001100110,
64'b1010101010101010101010101010101011000011001111001100001100111100,
64'b1100110000110011001100111100110011110000000011110000111111110000,
64'b0101101010100101101001010101101011000011001111001100001100111100,
64'b1111111100000000111111110000000001011010010110100101101001011010,
64'b0101101010100101101001010101101000000000000000000000000000000000,
64'b0011001111001100001100111100110010101010010101010101010110101010,
64'b1100110011001100110011001100110000111100001111000011110000111100,
64'b1100001111000011001111000011110010100101101001010101101001011010,
64'b0000111100001111111100001111000000000000111111111111111100000000,
64'b0000000000000000000000000000000000111100110000111100001100111100,
64'b1001011001101001011010011001011001010101101010100101010110101010,
64'b0101010110101010010101011010101010010110011010010110100110010110,
64'b1001011010010110100101101001011010010110100101101001011010010110,
64'b0101101001011010010110100101101011110000000011110000111111110000,
64'b1111111100000000111111110000000000000000111111111111111100000000,
64'b0110011001100110011001100110011001011010101001011010010101011010,
64'b0000111111110000000011111111000000110011110011000011001111001100,
64'b0000111111110000000011111111000010101010101010101010101010101010,
64'b1010010110100101010110100101101000110011001100111100110011001100,
64'b0101101010100101101001010101101010100101010110101010010101011010,
64'b0011001111001100001100111100110000110011110011000011001111001100,
64'b1111000000001111000011111111000001010101010101011010101010101010,
64'b1010101001010101010101011010101001011010101001011010010101011010,
64'b0000000000000000000000000000000010011001100110010110011001100110,
64'b1100110000110011001100111100110000111100110000111100001100111100,
64'b0101010101010101101010101010101001101001100101100110100110010110,
64'b1010010101011010101001010101101000000000111111111111111100000000,
64'b0000111111110000000011111111000001010101010101011010101010101010,
64'b0011110011000011110000110011110001100110100110011001100101100110,
64'b0101101001011010010110100101101001011010010110100101101001011010,
64'b0000000011111111111111110000000011001100110011001100110011001100,
64'b0011001111001100001100111100110011110000111100001111000011110000,
64'b0110011010011001100110010110011001100110100110011001100101100110,
64'b1010010110100101010110100101101000001111000011111111000011110000,
64'b0000000011111111111111110000000011001100110011001100110011001100,
64'b1001100110011001011001100110011001100110100110011001100101100110,
64'b1010101010101010101010101010101010010110100101101001011010010110,
64'b0000111100001111111100001111000001011010101001011010010101011010,
64'b0110011001100110011001100110011010010110011010010110100110010110,
64'b0110011010011001100110010110011011111111111111110000000000000000,
64'b0000000011111111111111110000000001100110011001100110011001100110,
64'b1111000000001111000011111111000001101001011010011001011010010110,
64'b1001100101100110100110010110011010011001011001101001100101100110,
64'b0101010101010101101010101010101001011010010110100101101001011010,
64'b1010010110100101010110100101101011111111000000001111111100000000,
64'b1100001111000011001111000011110011000011110000110011110000111100,
64'b1001100101100110100110010110011001010101101010100101010110101010,
64'b0101010101010101101010101010101001011010010110100101101001011010,
64'b1001011010010110100101101001011011000011110000110011110000111100,
64'b0110011001100110011001100110011001101001100101100110100110010110,
64'b1111111100000000111111110000000011001100001100110011001111001100,
64'b1001011010010110100101101001011010010110011010010110100110010110,
64'b1100001111000011001111000011110010101010101010101010101010101010,
64'b0101010101010101101010101010101010010110100101101001011010010110,
64'b1010101001010101010101011010101011000011001111001100001100111100,
64'b1001011010010110100101101001011010010110100101101001011010010110,
64'b1100110011001100110011001100110010011001011001101001100101100110,
64'b1001100101100110100110010110011011111111111111110000000000000000,
64'b1010010101011010101001010101101000001111111100000000111111110000,
64'b0110100101101001100101101001011010011001100110010110011001100110,
64'b1100110011001100110011001100110000110011110011000011001111001100,
64'b0110100110010110011010011001011000001111111100000000111111110000,
64'b0011110000111100001111000011110010010110011010010110100110010110,
64'b1111111111111111000000000000000000001111000011111111000011110000,
64'b1100001100111100110000110011110010010110011010010110100110010110,
64'b0000111111110000000011111111000001100110011001100110011001100110,
64'b0110011001100110011001100110011011000011001111001100001100111100,
64'b1001100110011001011001100110011011110000000011110000111111110000,
64'b0110100110010110011010011001011011000011001111001100001100111100,
64'b1010010110100101010110100101101011111111111111110000000000000000,
64'b1100001111000011001111000011110011001100110011001100110011001100,
64'b1010101001010101010101011010101010011001011001101001100101100110,
64'b0011110011000011110000110011110010100101010110101010010101011010,
64'b1010010101011010101001010101101000111100110000111100001100111100,
64'b0000111111110000000011111111000000001111111100000000111111110000,
64'b0101010110101010010101011010101000111100110000111100001100111100,
64'b0000111100001111111100001111000001101001100101100110100110010110,
64'b1111000000001111000011111111000010101010010101010101010110101010,
64'b0110011010011001100110010110011001010101101010100101010110101010,
64'b0011001111001100001100111100110001101001011010011001011010010110,
64'b0101010101010101101010101010101001100110011001100110011001100110,
64'b1100001100111100110000110011110001011010010110100101101001011010,
64'b0011110011000011110000110011110000000000000000000000000000000000,
64'b0110011010011001100110010110011001011010010110100101101001011010,
64'b0011001111001100001100111100110011000011110000110011110000111100,
64'b0110011001100110011001100110011011001100001100110011001111001100,
64'b1100001111000011001111000011110011110000000011110000111111110000,
64'b0000111100001111111100001111000010101010010101010101010110101010,
64'b0110011010011001100110010110011011110000000011110000111111110000,
64'b1111000000001111000011111111000010010110011010010110100110010110,
64'b0101101001011010010110100101101000110011001100111100110011001100,
64'b0000111111110000000011111111000010011001100110010110011001100110,
64'b1001011001101001011010011001011011000011001111001100001100111100,
64'b1001100110011001011001100110011010010110100101101001011010010110,
64'b0110011001100110011001100110011000110011110011000011001111001100,
64'b0101010110101010010101011010101000000000000000000000000000000000,
64'b1010101010101010101010101010101000110011110011000011001111001100,
64'b0000111111110000000011111111000000001111111100000000111111110000,
64'b0000000011111111111111110000000010100101101001010101101001011010,
64'b1010101010101010101010101010101010101010010101010101010110101010,
64'b0101101001011010010110100101101010011001100110010110011001100110,
64'b0011110011000011110000110011110010101010010101010101010110101010,
64'b1010010101011010101001010101101010010110011010010110100110010110,
64'b0110100101101001100101101001011001011010010110100101101001011010,
64'b0110011001100110011001100110011010010110100101101001011010010110,
64'b0000111100001111111100001111000001011010101001011010010101011010,
64'b1100001111000011001111000011110011000011001111001100001100111100,
64'b0101010110101010010101011010101011110000111100001111000011110000,
64'b0011001100110011110011001100110010101010101010101010101010101010,
64'b1100110011001100110011001100110000001111000011111111000011110000,
64'b0000000011111111111111110000000000000000111111111111111100000000,
64'b1111111111111111000000000000000000110011110011000011001111001100,
64'b0110011001100110011001100110011010011001100110010110011001100110,
64'b0011001111001100001100111100110010010110100101101001011010010110,
64'b1111000000001111000011111111000010011001100110010110011001100110,
64'b0110011010011001100110010110011010010110011010010110100110010110,
64'b1100001100111100110000110011110010011001011001101001100101100110,
64'b1001011010010110100101101001011011000011001111001100001100111100,
64'b1111111100000000111111110000000011001100001100110011001111001100,
64'b1010010101011010101001010101101001011010101001011010010101011010,
64'b0110011001100110011001100110011011111111000000001111111100000000,
64'b0101010101010101101010101010101011001100110011001100110011001100,
64'b1001100110011001011001100110011011111111000000001111111100000000,
64'b0101010110101010010101011010101001010101010101011010101010101010,
64'b1001011001101001011010011001011010100101101001010101101001011010,
64'b0011001111001100001100111100110000111100001111000011110000111100,
64'b0000000011111111111111110000000001101001100101100110100110010110,
64'b0101010101010101101010101010101000111100001111000011110000111100,
64'b0110011001100110011001100110011010010110011010010110100110010110,
64'b1010101010101010101010101010101001101001011010011001011010010110,
64'b1010010110100101010110100101101011110000000011110000111111110000,
64'b1100110000110011001100111100110000001111000011111111000011110000,
64'b1001100101100110100110010110011001100110100110011001100101100110,
64'b1111111100000000111111110000000010101010101010101010101010101010,
64'b1100001111000011001111000011110001011010010110100101101001011010,
64'b0101010101010101101010101010101011111111111111110000000000000000,
64'b0011001111001100001100111100110011001100110011001100110011001100,
64'b0000000000000000000000000000000010011001011001101001100101100110,
64'b0000000011111111111111110000000010100101010110101010010101011010,
64'b1111000000001111000011111111000000111100110000111100001100111100,
64'b0011001111001100001100111100110000001111111100000000111111110000,
64'b1001100110011001011001100110011000111100110000111100001100111100,
64'b0011110011000011110000110011110001101001100101100110100110010110,
64'b0101010101010101101010101010101010101010010101010101010110101010,
64'b1001011001101001011010011001011001010101101010100101010110101010,
64'b0011110000111100001111000011110001101001011010011001011010010110,
64'b1100001100111100110000110011110001100110011001100110011001100110,
64'b1010010101011010101001010101101000111100110000111100001100111100,
64'b0110011001100110011001100110011011000011110000110011110000111100,
64'b1010010110100101010110100101101011110000000011110000111111110000,
64'b0000000000000000000000000000000011111111000000001111111100000000,
64'b1111111111111111000000000000000001101001011010011001011010010110,
64'b1010101001010101010101011010101011111111111111110000000000000000,
64'b1010010110100101010110100101101011111111111111110000000000000000,
64'b0011110000111100001111000011110011111111000000001111111100000000,
64'b0101101010100101101001010101101001100110011001100110011001100110,
64'b0110011001100110011001100110011001010101101010100101010110101010,
64'b1001011001101001011010011001011010101010010101010101010110101010,
64'b1010010101011010101001010101101010010110011010010110100110010110,
64'b0000111111110000000011111111000001010101101010100101010110101010,
64'b1100001100111100110000110011110001010101101010100101010110101010,
64'b1111111111111111000000000000000001100110100110011001100101100110,
64'b1001100110011001011001100110011000000000000000000000000000000000,
64'b1001011001101001011010011001011001101001100101100110100110010110,
64'b1010010101011010101001010101101001100110011001100110011001100110,
64'b1001011001101001011010011001011010100101010110101010010101011010,
64'b1100110011001100110011001100110011111111000000001111111100000000,
64'b1010101001010101010101011010101001011010010110100101101001011010,
64'b0011110000111100001111000011110011001100001100110011001111001100,
64'b1111000000001111000011111111000001010101101010100101010110101010,
64'b0000111100001111111100001111000000000000111111111111111100000000,
64'b0011001111001100001100111100110011000011001111001100001100111100,
64'b0011110000111100001111000011110010100101010110101010010101011010,
64'b1111111100000000111111110000000010011001100110010110011001100110,
64'b1100001111000011001111000011110011000011110000110011110000111100,
64'b0011110011000011110000110011110010101010101010101010101010101010,
64'b1010101010101010101010101010101000111100110000111100001100111100,
64'b1100001111000011001111000011110000111100001111000011110000111100,
64'b0011001100110011110011001100110011001100001100110011001111001100,
64'b0000111111110000000011111111000011111111111111110000000000000000,
64'b0011110000111100001111000011110000110011110011000011001111001100,
64'b0101010101010101101010101010101000001111000011111111000011110000,
64'b0110011001100110011001100110011010011001100110010110011001100110,
64'b0110011001100110011001100110011011111111111111110000000000000000,
64'b1111000011110000111100001111000001011010101001011010010101011010,
64'b1100110011001100110011001100110000110011110011000011001111001100,
64'b1111111111111111000000000000000010010110100101101001011010010110,
64'b0000111111110000000011111111000010100101010110101010010101011010,
64'b0101101010100101101001010101101001100110011001100110011001100110,
64'b0110011001100110011001100110011011110000000011110000111111110000,
64'b0000111111110000000011111111000010100101010110101010010101011010,
64'b0101101001011010010110100101101000001111000011111111000011110000,
64'b1010101001010101010101011010101010101010101010101010101010101010,
64'b0000111111110000000011111111000010100101101001010101101001011010,
64'b1100110011001100110011001100110011111111000000001111111100000000,
64'b1001011010010110100101101001011010010110100101101001011010010110,
64'b0011110000111100001111000011110010101010101010101010101010101010,
64'b1111111100000000111111110000000001100110100110011001100101100110,
64'b1111000011110000111100001111000001011010010110100101101001011010,
64'b1010010110100101010110100101101001100110100110011001100101100110,
64'b0110100110010110011010011001011000001111111100000000111111110000,
64'b0110011001100110011001100110011010010110011010010110100110010110,
64'b1010101001010101010101011010101000111100001111000011110000111100,
64'b1010010110100101010110100101101011000011110000110011110000111100,
64'b0011110000111100001111000011110011110000111100001111000011110000,
64'b0110011010011001100110010110011000110011110011000011001111001100,
64'b1010010101011010101001010101101000111100110000111100001100111100,
64'b0000000011111111111111110000000010100101010110101010010101011010,
64'b1010010110100101010110100101101010100101101001010101101001011010,
64'b0011110000111100001111000011110011111111000000001111111100000000,
64'b1010101010101010101010101010101010010110100101101001011010010110,
64'b0011110000111100001111000011110001011010010110100101101001011010,
64'b0011110011000011110000110011110011000011110000110011110000111100,
64'b0101010110101010010101011010101010101010010101010101010110101010,
64'b1001011001101001011010011001011000111100110000111100001100111100,
64'b0000111111110000000011111111000010100101010110101010010101011010,
64'b0011110000111100001111000011110000001111111100000000111111110000,
64'b1010101010101010101010101010101001010101101010100101010110101010,
64'b1001011001101001011010011001011000001111000011111111000011110000,
64'b0110100110010110011010011001011011110000000011110000111111110000,
64'b0000111111110000000011111111000001100110100110011001100101100110,
64'b1111111111111111000000000000000000110011110011000011001111001100,
64'b1001011010010110100101101001011001010101010101011010101010101010,
64'b1001100110011001011001100110011011000011001111001100001100111100,
64'b1100110011001100110011001100110000110011110011000011001111001100,
64'b1111111100000000111111110000000010100101010110101010010101011010,
64'b0101101001011010010110100101101010011001100110010110011001100110,
64'b1001011010010110100101101001011001011010101001011010010101011010,
64'b1001011010010110100101101001011001100110100110011001100101100110,
64'b1010101010101010101010101010101000000000111111111111111100000000,
64'b1100001100111100110000110011110000110011001100111100110011001100,
64'b0110100101101001100101101001011011111111000000001111111100000000,
64'b1001100101100110100110010110011010101010010101010101010110101010,
64'b1111000011110000111100001111000001101001011010011001011010010110,
64'b0110011010011001100110010110011010100101101001010101101001011010,
64'b0101101001011010010110100101101011001100110011001100110011001100,
64'b0110100101101001100101101001011001011010101001011010010101011010,
64'b1001100101100110100110010110011011110000111100001111000011110000,
64'b1111111111111111000000000000000011001100001100110011001111001100,
64'b0011001111001100001100111100110000111100001111000011110000111100,
64'b1100001100111100110000110011110001100110100110011001100101100110,
64'b1100001100111100110000110011110001101001011010011001011010010110,
64'b1100110011001100110011001100110001010101010101011010101010101010,
64'b1111000000001111000011111111000001011010010110100101101001011010,
64'b1100001100111100110000110011110001010101010101011010101010101010,
64'b0110100101101001100101101001011000110011001100111100110011001100,
64'b1111111100000000111111110000000001101001100101100110100110010110,
64'b1100001111000011001111000011110010011001011001101001100101100110,
64'b1001100101100110100110010110011001011010010110100101101001011010,
64'b1100001100111100110000110011110011001100001100110011001111001100,
64'b1001011010010110100101101001011001010101101010100101010110101010,
64'b1010101010101010101010101010101010100101101001010101101001011010,
64'b1010010110100101010110100101101010100101010110101010010101011010,
64'b1111000000001111000011111111000011000011110000110011110000111100,
64'b1111000000001111000011111111000001101001100101100110100110010110,
64'b1111000011110000111100001111000001100110011001100110011001100110,
64'b0000000011111111111111110000000010011001011001101001100101100110,
64'b0101101010100101101001010101101011001100110011001100110011001100,
64'b1100001100111100110000110011110001011010010110100101101001011010,
64'b0101010101010101101010101010101010010110011010010110100110010110,
64'b0000111111110000000011111111000011000011110000110011110000111100,
64'b0110100101101001100101101001011000110011110011000011001111001100,
64'b1111000000001111000011111111000000001111000011111111000011110000,
64'b1100001100111100110000110011110001100110011001100110011001100110,
64'b1100110011001100110011001100110000110011110011000011001111001100,
64'b0011001111001100001100111100110001100110100110011001100101100110,
64'b1010101001010101010101011010101000001111111100000000111111110000,
64'b1010101001010101010101011010101010010110011010010110100110010110,
64'b0101010110101010010101011010101000111100001111000011110000111100,
64'b1111111111111111000000000000000011000011110000110011110000111100,
64'b0110011010011001100110010110011011110000111100001111000011110000,
64'b0101101010100101101001010101101000110011110011000011001111001100,
64'b1100110011001100110011001100110000111100110000111100001100111100,
64'b1010101001010101010101011010101010100101010110101010010101011010,
64'b1100001100111100110000110011110010100101101001010101101001011010,
64'b1010101001010101010101011010101011111111000000001111111100000000,
64'b1010010101011010101001010101101010010110100101101001011010010110,
64'b0000111100001111111100001111000010010110011010010110100110010110,
64'b0000111100001111111100001111000000110011001100111100110011001100,
64'b0110011001100110011001100110011000000000111111111111111100000000,
64'b0110100101101001100101101001011001010101101010100101010110101010,
64'b1010101001010101010101011010101011110000000011110000111111110000,
64'b1100001100111100110000110011110010101010010101010101010110101010,
64'b0110011010011001100110010110011000110011001100111100110011001100,
64'b0110100101101001100101101001011010011001011001101001100101100110,
64'b1100110000110011001100111100110010100101101001010101101001011010,
64'b0000111111110000000011111111000011111111111111110000000000000000,
64'b1010101001010101010101011010101001011010101001011010010101011010,
64'b1100110011001100110011001100110011111111111111110000000000000000,
64'b1010101010101010101010101010101001010101101010100101010110101010,
64'b0101101010100101101001010101101000111100110000111100001100111100,
64'b0101101010100101101001010101101001011010010110100101101001011010,
64'b1111000011110000111100001111000001010101010101011010101010101010,
64'b1010101001010101010101011010101010011001100110010110011001100110,
64'b0011001111001100001100111100110000000000111111111111111100000000,
64'b1001100110011001011001100110011010011001100110010110011001100110,
64'b1010010101011010101001010101101001011010010110100101101001011010,
64'b0000000011111111111111110000000001101001011010011001011010010110,
64'b0110100110010110011010011001011000110011110011000011001111001100,
64'b1010010110100101010110100101101010101010101010101010101010101010,
64'b1001100101100110100110010110011001100110100110011001100101100110,
64'b1001011010010110100101101001011010101010101010101010101010101010,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b1100001100111100110000110011110001011010101001011010010101011010,
64'b0110100110010110011010011001011010011001011001101001100101100110,
64'b0011001111001100001100111100110011001100110011001100110011001100,
64'b0101101001011010010110100101101010010110100101101001011010010110,
64'b0000111111110000000011111111000001010101010101011010101010101010,
64'b1111111100000000111111110000000010010110100101101001011010010110,
64'b0000000000000000000000000000000010011001011001101001100101100110,
64'b1001011010010110100101101001011011000011001111001100001100111100,
64'b0101101001011010010110100101101010100101101001010101101001011010,
64'b0011110000111100001111000011110011001100110011001100110011001100,
64'b1100001100111100110000110011110011000011110000110011110000111100,
64'b0000111111110000000011111111000001100110011001100110011001100110,
64'b1001011010010110100101101001011000111100001111000011110000111100,
64'b0101101010100101101001010101101011001100001100110011001111001100,
64'b0011110011000011110000110011110001101001011010011001011010010110,
64'b0000111100001111111100001111000011110000111100001111000011110000,
64'b0011001111001100001100111100110011000011001111001100001100111100,
64'b0000000011111111111111110000000011001100110011001100110011001100,
64'b1111111111111111000000000000000001101001100101100110100110010110,
64'b0000000000000000000000000000000011000011110000110011110000111100,
64'b1100001100111100110000110011110011110000000011110000111111110000,
64'b0011001111001100001100111100110000110011110011000011001111001100,
64'b0000111111110000000011111111000001011010010110100101101001011010,
64'b1111000000001111000011111111000000001111111100000000111111110000,
64'b0000000011111111111111110000000010010110100101101001011010010110,
64'b1100001100111100110000110011110000001111111100000000111111110000,
64'b1100001100111100110000110011110010100101101001010101101001011010,
64'b0101010110101010010101011010101001101001100101100110100110010110,
64'b0011001111001100001100111100110001010101101010100101010110101010,
64'b1100110011001100110011001100110011110000000011110000111111110000,
64'b0101010110101010010101011010101011110000111100001111000011110000,
64'b0110100110010110011010011001011000111100110000111100001100111100,
64'b1100110000110011001100111100110000001111111100000000111111110000,
64'b1001100101100110100110010110011010101010010101010101010110101010,
64'b1100001100111100110000110011110010100101101001010101101001011010,
64'b0000111100001111111100001111000000110011110011000011001111001100,
64'b1010101010101010101010101010101000000000111111111111111100000000,
64'b1001100110011001011001100110011011000011001111001100001100111100,
64'b0000111111110000000011111111000011111111000000001111111100000000,
64'b0101010110101010010101011010101000110011110011000011001111001100,
64'b0011110000111100001111000011110010010110011010010110100110010110,
64'b0110100101101001100101101001011000110011001100111100110011001100,
64'b1001100110011001011001100110011000000000111111111111111100000000,
64'b1001100101100110100110010110011001010101101010100101010110101010,
64'b1111111111111111000000000000000011110000000011110000111111110000,
64'b0110100110010110011010011001011010101010010101010101010110101010,
64'b0000000000000000000000000000000000110011001100111100110011001100,
64'b0011110000111100001111000011110010011001011001101001100101100110,
64'b1111000011110000111100001111000010100101101001010101101001011010,
64'b1100110000110011001100111100110011111111111111110000000000000000,
64'b1111000011110000111100001111000001011010101001011010010101011010,
64'b1111111100000000111111110000000000000000000000000000000000000000,
64'b1001100110011001011001100110011000000000000000000000000000000000,
64'b0000111111110000000011111111000000110011110011000011001111001100,
64'b1100001100111100110000110011110000111100001111000011110000111100,
64'b1001011010010110100101101001011000111100001111000011110000111100,
64'b0110100101101001100101101001011000110011110011000011001111001100,
64'b0000000000000000000000000000000011000011110000110011110000111100,
64'b1001011001101001011010011001011011111111000000001111111100000000,
64'b0000000000000000000000000000000000110011001100111100110011001100,
64'b0000111111110000000011111111000010100101010110101010010101011010,
64'b1111111100000000111111110000000000111100001111000011110000111100,
64'b0000111100001111111100001111000000000000111111111111111100000000,
64'b0101010110101010010101011010101010101010010101010101010110101010,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1001100110011001011001100110011010100101101001010101101001011010,
64'b1010010101011010101001010101101000000000000000000000000000000000,
64'b1001011001101001011010011001011001101001100101100110100110010110,
64'b1010101001010101010101011010101001100110100110011001100101100110,
64'b0110100101101001100101101001011010100101010110101010010101011010,
64'b0110100110010110011010011001011011001100110011001100110011001100,
64'b0101101001011010010110100101101000110011110011000011001111001100,
64'b1100001111000011001111000011110010011001100110010110011001100110,
64'b1100110011001100110011001100110010101010101010101010101010101010,
64'b1111000000001111000011111111000000000000000000000000000000000000,
64'b0101010101010101101010101010101001010101101010100101010110101010,
64'b0101010101010101101010101010101001010101010101011010101010101010,
64'b1010101010101010101010101010101000000000000000000000000000000000,
64'b0011001100110011110011001100110010011001011001101001100101100110,
64'b0110100110010110011010011001011010101010101010101010101010101010,
64'b0101101010100101101001010101101000111100110000111100001100111100,
64'b1111000011110000111100001111000011000011110000110011110000111100,
64'b1100001111000011001111000011110001100110100110011001100101100110,
64'b0101010101010101101010101010101011110000111100001111000011110000,
64'b0101010101010101101010101010101000001111000011111111000011110000,
64'b0110011010011001100110010110011000111100001111000011110000111100,
64'b1001011001101001011010011001011001100110011001100110011001100110,
64'b0000111100001111111100001111000000000000000000000000000000000000,
64'b1100110000110011001100111100110000110011001100111100110011001100,
64'b1010101010101010101010101010101011001100110011001100110011001100,
64'b1100110011001100110011001100110010101010101010101010101010101010,
64'b1111000011110000111100001111000001101001011010011001011010010110,
64'b1001011001101001011010011001011011001100110011001100110011001100,
64'b1100110000110011001100111100110011110000000011110000111111110000,
64'b0101010110101010010101011010101010100101010110101010010101011010,
64'b0000111111110000000011111111000001101001011010011001011010010110,
64'b0110011001100110011001100110011001010101101010100101010110101010,
64'b0110011001100110011001100110011011111111000000001111111100000000,
64'b0110100101101001100101101001011010100101010110101010010101011010,
64'b1001011001101001011010011001011000111100001111000011110000111100,
64'b0101010110101010010101011010101000000000000000000000000000000000,
64'b1010010110100101010110100101101011110000111100001111000011110000,
64'b0110011001100110011001100110011001011010010110100101101001011010,
64'b1111000011110000111100001111000011001100110011001100110011001100,
64'b1111000000001111000011111111000011001100001100110011001111001100,
64'b0011001111001100001100111100110001010101010101011010101010101010,
64'b1100001111000011001111000011110001100110100110011001100101100110,
64'b1111000011110000111100001111000000001111111100000000111111110000,
64'b1010101010101010101010101010101001101001011010011001011010010110,
64'b1111111100000000111111110000000001011010101001011010010101011010,
64'b0101101010100101101001010101101010011001011001101001100101100110,
64'b1010101001010101010101011010101010100101010110101010010101011010,
64'b0101101001011010010110100101101011000011110000110011110000111100,
64'b1001011001101001011010011001011000001111111100000000111111110000,
64'b1001100110011001011001100110011001010101010101011010101010101010,
64'b0101101001011010010110100101101011111111000000001111111100000000,
64'b0101010110101010010101011010101001011010010110100101101001011010,
64'b0000111111110000000011111111000000001111000011111111000011110000,
64'b1010101010101010101010101010101001100110011001100110011001100110,
64'b0110100110010110011010011001011001101001011010011001011010010110,
64'b0011110011000011110000110011110010101010010101010101010110101010,
64'b0110011010011001100110010110011011000011001111001100001100111100,
64'b0011110011000011110000110011110001100110100110011001100101100110,
64'b1010101010101010101010101010101001101001011010011001011010010110,
64'b1111000011110000111100001111000011001100001100110011001111001100,
64'b0101010101010101101010101010101000001111111100000000111111110000,
64'b0011001100110011110011001100110010101010010101010101010110101010,
64'b0011110011000011110000110011110011001100110011001100110011001100,
64'b0101010110101010010101011010101001010101010101011010101010101010,
64'b0110011001100110011001100110011000110011110011000011001111001100,
64'b0000111111110000000011111111000001010101101010100101010110101010,
64'b1100001111000011001111000011110010010110100101101001011010010110,
64'b0101101010100101101001010101101011000011001111001100001100111100,
64'b1001100101100110100110010110011010011001100110010110011001100110,
64'b1100001100111100110000110011110001011010101001011010010101011010,
64'b1001100110011001011001100110011011000011110000110011110000111100,
64'b0000000011111111111111110000000001101001100101100110100110010110,
64'b1001011001101001011010011001011010100101101001010101101001011010,
64'b0000000011111111111111110000000010101010010101010101010110101010,
64'b0101010110101010010101011010101000110011001100111100110011001100,
64'b1111000011110000111100001111000001011010010110100101101001011010,
64'b0101010101010101101010101010101011001100110011001100110011001100,
64'b1001011010010110100101101001011001011010010110100101101001011010,
64'b1010101001010101010101011010101000110011001100111100110011001100,
64'b0000111111110000000011111111000011000011001111001100001100111100,
64'b0110011010011001100110010110011011110000000011110000111111110000,
64'b0110100101101001100101101001011000111100001111000011110000111100,
64'b1111000000001111000011111111000001100110100110011001100101100110,
64'b0011110000111100001111000011110010100101010110101010010101011010,
64'b0101010101010101101010101010101010010110011010010110100110010110,
64'b1001011001101001011010011001011000110011110011000011001111001100,
64'b0101010101010101101010101010101010011001100110010110011001100110,
64'b1001100110011001011001100110011001011010010110100101101001011010,
64'b1111111100000000111111110000000010011001011001101001100101100110,
64'b1100110011001100110011001100110011110000111100001111000011110000,
64'b0110100110010110011010011001011000110011110011000011001111001100,
64'b0011001100110011110011001100110001011010010110100101101001011010,
64'b1010101001010101010101011010101001011010101001011010010101011010,
64'b1100001111000011001111000011110000000000111111111111111100000000,
64'b0110100110010110011010011001011010100101010110101010010101011010,
64'b1010101001010101010101011010101011000011110000110011110000111100,
64'b1010010101011010101001010101101001100110100110011001100101100110,
64'b1100110011001100110011001100110000111100110000111100001100111100,
64'b1001011001101001011010011001011010100101101001010101101001011010,
64'b0110011001100110011001100110011000111100001111000011110000111100,
64'b1001011010010110100101101001011010011001011001101001100101100110,
64'b0101010101010101101010101010101011000011110000110011110000111100,
64'b1111000011110000111100001111000011111111000000001111111100000000,
64'b1100001100111100110000110011110011110000111100001111000011110000,
64'b0101101001011010010110100101101000110011110011000011001111001100,
64'b1001100110011001011001100110011011001100001100110011001111001100,
64'b1010010101011010101001010101101001010101010101011010101010101010,
64'b1001011001101001011010011001011001100110100110011001100101100110,
64'b0011001100110011110011001100110000001111111100000000111111110000,
64'b0110011010011001100110010110011001101001011010011001011010010110,
64'b1111000011110000111100001111000001011010101001011010010101011010,
64'b0011110011000011110000110011110010011001011001101001100101100110,
64'b1001011010010110100101101001011010100101010110101010010101011010,
64'b1100001100111100110000110011110011000011110000110011110000111100,
64'b1100110011001100110011001100110000001111111100000000111111110000,
64'b0101010110101010010101011010101001010101010101011010101010101010,
64'b0000111111110000000011111111000011111111000000001111111100000000,
64'b1010010110100101010110100101101011001100110011001100110011001100,
64'b1100110000110011001100111100110011000011110000110011110000111100,
64'b0000111111110000000011111111000000000000111111111111111100000000,
64'b1001100101100110100110010110011001010101101010100101010110101010,
64'b0000000000000000000000000000000001011010101001011010010101011010,
64'b1001011001101001011010011001011011111111111111110000000000000000,
64'b0101101010100101101001010101101000110011001100111100110011001100,
64'b1010101010101010101010101010101001100110100110011001100101100110,
64'b1010101010101010101010101010101011111111111111110000000000000000,
64'b1100001111000011001111000011110001010101010101011010101010101010,
64'b1100110000110011001100111100110001101001100101100110100110010110,
64'b0101010110101010010101011010101000110011001100111100110011001100,
64'b1001011010010110100101101001011011110000111100001111000011110000,
64'b1001011001101001011010011001011001011010010110100101101001011010,
64'b0110100110010110011010011001011000001111111100000000111111110000,
64'b1010010110100101010110100101101001010101010101011010101010101010,
64'b0101101010100101101001010101101010011001100110010110011001100110,
64'b0000000000000000000000000000000011001100001100110011001111001100,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b0011110000111100001111000011110001011010010110100101101001011010,
64'b1100110011001100110011001100110001101001011010011001011010010110,
64'b0110011001100110011001100110011010101010101010101010101010101010,
64'b1100110000110011001100111100110001100110011001100110011001100110,
64'b0110100110010110011010011001011010010110011010010110100110010110,
64'b1100110000110011001100111100110011110000111100001111000011110000,
64'b0101010110101010010101011010101001010101101010100101010110101010,
64'b1001100101100110100110010110011000110011110011000011001111001100,
64'b0101101001011010010110100101101000000000111111111111111100000000,
64'b0011110000111100001111000011110011001100110011001100110011001100,
64'b1111111111111111000000000000000010010110100101101001011010010110,
64'b1010101010101010101010101010101010100101101001010101101001011010,
64'b0101101010100101101001010101101001100110011001100110011001100110,
64'b0101010101010101101010101010101000110011110011000011001111001100,
64'b0101101001011010010110100101101011000011001111001100001100111100,
64'b1001011010010110100101101001011001100110011001100110011001100110,
64'b1100110011001100110011001100110000111100001111000011110000111100,
64'b0101101001011010010110100101101000111100110000111100001100111100,
64'b0101101010100101101001010101101001010101101010100101010110101010,
64'b1111000011110000111100001111000011001100110011001100110011001100,
64'b1100001111000011001111000011110000001111000011111111000011110000,
64'b0011001111001100001100111100110011111111111111110000000000000000,
64'b0000111111110000000011111111000001011010010110100101101001011010,
64'b0000000000000000000000000000000011000011001111001100001100111100,
64'b0110011001100110011001100110011000110011110011000011001111001100,
64'b1100110000110011001100111100110010010110100101101001011010010110,
64'b0110011001100110011001100110011000001111000011111111000011110000,
64'b1001100101100110100110010110011011110000000011110000111111110000,
64'b1100001100111100110000110011110000111100001111000011110000111100,
64'b1111000011110000111100001111000000001111111100000000111111110000,
64'b0011001111001100001100111100110011110000000011110000111111110000,
64'b1100110000110011001100111100110010011001100110010110011001100110,
64'b0101010110101010010101011010101011110000111100001111000011110000,
64'b0000000011111111111111110000000001010101101010100101010110101010,
64'b0110100110010110011010011001011010101010101010101010101010101010,
64'b0000111100001111111100001111000010011001011001101001100101100110,
64'b1001100101100110100110010110011011110000000011110000111111110000,
64'b0011110000111100001111000011110000001111000011111111000011110000,
64'b1001100101100110100110010110011011000011001111001100001100111100,
64'b1100110000110011001100111100110011111111000000001111111100000000,
64'b0110100101101001100101101001011010101010010101010101010110101010,
64'b0101101010100101101001010101101010100101010110101010010101011010,
64'b0011110011000011110000110011110000000000111111111111111100000000,
64'b1100001100111100110000110011110000000000111111111111111100000000,
64'b0101101010100101101001010101101010010110100101101001011010010110,
64'b1111000011110000111100001111000001010101101010100101010110101010,
64'b1111000011110000111100001111000010011001100110010110011001100110,
64'b0101101001011010010110100101101011001100110011001100110011001100,
64'b1111000011110000111100001111000011000011110000110011110000111100,
64'b1111000000001111000011111111000000000000111111111111111100000000,
64'b0000111111110000000011111111000001010101101010100101010110101010,
64'b0101010110101010010101011010101001011010101001011010010101011010,
64'b0101010110101010010101011010101011111111111111110000000000000000,
64'b1100001100111100110000110011110000110011001100111100110011001100,
64'b1100110000110011001100111100110001100110100110011001100101100110,
64'b1001100101100110100110010110011011111111111111110000000000000000,
64'b1001011010010110100101101001011001010101010101011010101010101010,
64'b1001100110011001011001100110011001101001100101100110100110010110,
64'b1100001100111100110000110011110011001100110011001100110011001100,
64'b0101010110101010010101011010101010011001100110010110011001100110,
64'b0011001111001100001100111100110010010110011010010110100110010110,
64'b1111111100000000111111110000000000000000000000000000000000000000,
64'b0000000011111111111111110000000011001100001100110011001111001100,
64'b1010101001010101010101011010101010011001100110010110011001100110,
64'b0011001100110011110011001100110001011010010110100101101001011010,
64'b0011001100110011110011001100110011110000000011110000111111110000,
64'b1111000000001111000011111111000011110000111100001111000011110000,
64'b0000111100001111111100001111000011000011110000110011110000111100,
64'b0110100101101001100101101001011001101001011010011001011010010110,
64'b1100001100111100110000110011110010101010010101010101010110101010,
64'b0011110000111100001111000011110011000011110000110011110000111100,
64'b1010010101011010101001010101101001100110011001100110011001100110,
64'b1001011010010110100101101001011010011001100110010110011001100110,
64'b1100001100111100110000110011110001011010010110100101101001011010,
64'b1111000000001111000011111111000010100101010110101010010101011010,
64'b0110011010011001100110010110011010010110011010010110100110010110,
64'b1001100110011001011001100110011010010110100101101001011010010110,
64'b1100110000110011001100111100110000001111000011111111000011110000,
64'b0000000011111111111111110000000001011010010110100101101001011010,
64'b0000000011111111111111110000000011111111000000001111111100000000,
64'b1111111100000000111111110000000010100101010110101010010101011010,
64'b1010101001010101010101011010101010101010010101010101010110101010,
64'b1001011010010110100101101001011001010101101010100101010110101010,
64'b0101101001011010010110100101101011110000111100001111000011110000,
64'b1010010101011010101001010101101000000000000000000000000000000000,
64'b0110011010011001100110010110011000111100001111000011110000111100,
64'b0011110000111100001111000011110010011001011001101001100101100110,
64'b0000111100001111111100001111000011001100001100110011001111001100,
64'b1111000000001111000011111111000000111100110000111100001100111100,
64'b1001011010010110100101101001011001101001100101100110100110010110,
64'b0011001111001100001100111100110011111111000000001111111100000000,
64'b0000111111110000000011111111000010011001011001101001100101100110,
64'b1111111111111111000000000000000011111111111111110000000000000000,
64'b1111111111111111000000000000000011001100001100110011001111001100,
64'b1111000011110000111100001111000000110011001100111100110011001100,
64'b1010010110100101010110100101101010011001100110010110011001100110,
64'b0110011001100110011001100110011011111111000000001111111100000000,
64'b1010010101011010101001010101101000000000000000000000000000000000,
64'b1100001111000011001111000011110000001111111100000000111111110000,
64'b1010010101011010101001010101101011000011110000110011110000111100,
64'b1111111100000000111111110000000000001111000011111111000011110000,
64'b1010101001010101010101011010101001011010101001011010010101011010,
64'b0110100110010110011010011001011010010110011010010110100110010110,
64'b0000111100001111111100001111000011111111111111110000000000000000,
64'b0000000011111111111111110000000011000011110000110011110000111100,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1010101010101010101010101010101010100101101001010101101001011010,
64'b0101010110101010010101011010101001011010010110100101101001011010,
64'b0011001111001100001100111100110010010110100101101001011010010110,
64'b1001011010010110100101101001011001010101010101011010101010101010,
64'b0011001111001100001100111100110000000000000000000000000000000000,
64'b1010101001010101010101011010101010100101010110101010010101011010,
64'b1010101010101010101010101010101011000011110000110011110000111100,
64'b1111000000001111000011111111000001011010010110100101101001011010,
64'b1010101001010101010101011010101011111111111111110000000000000000,
64'b1001011001101001011010011001011010010110011010010110100110010110,
64'b0110100101101001100101101001011000111100110000111100001100111100,
64'b0000111111110000000011111111000011111111111111110000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0110011001100110011001100110011010011001011001101001100101100110,
64'b1111000011110000111100001111000001011010101001011010010101011010,
64'b1100001100111100110000110011110000001111000011111111000011110000,
64'b1001011010010110100101101001011010011001011001101001100101100110,
64'b0110011001100110011001100110011000111100001111000011110000111100,
64'b0011110000111100001111000011110011001100001100110011001111001100,
64'b1010101001010101010101011010101000001111111100000000111111110000,
64'b0000111100001111111100001111000010011001011001101001100101100110,
64'b0000000011111111111111110000000000000000000000000000000000000000,
64'b1001011001101001011010011001011010010110011010010110100110010110,
64'b1111111111111111000000000000000001011010101001011010010101011010,
64'b1111000011110000111100001111000010101010101010101010101010101010,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b1001011010010110100101101001011011000011110000110011110000111100,
64'b0011110011000011110000110011110011001100001100110011001111001100,
64'b0011110000111100001111000011110001010101101010100101010110101010,
64'b1001011010010110100101101001011001101001011010011001011010010110,
64'b1010101010101010101010101010101000001111111100000000111111110000,
64'b1010101001010101010101011010101010100101101001010101101001011010,
64'b1111111100000000111111110000000010101010010101010101010110101010,
64'b0101101001011010010110100101101011000011110000110011110000111100,
64'b1100110000110011001100111100110000000000000000000000000000000000,
64'b1001011001101001011010011001011000111100110000111100001100111100,
64'b0011110011000011110000110011110001100110100110011001100101100110,
64'b0000111100001111111100001111000001100110011001100110011001100110,
64'b0110011001100110011001100110011011001100110011001100110011001100,
64'b0110100110010110011010011001011000001111111100000000111111110000,
64'b0011001111001100001100111100110010100101101001010101101001011010,
64'b0110100101101001100101101001011010011001100110010110011001100110,
64'b1001011010010110100101101001011011000011001111001100001100111100,
64'b0101101001011010010110100101101001010101101010100101010110101010,
64'b0011001100110011110011001100110000110011110011000011001111001100,
64'b0101010101010101101010101010101010011001100110010110011001100110,
64'b0011001111001100001100111100110010100101010110101010010101011010,
64'b0000111100001111111100001111000010101010101010101010101010101010,
64'b1001011001101001011010011001011011110000000011110000111111110000,
64'b0101101010100101101001010101101001101001011010011001011010010110,
64'b0101010110101010010101011010101010010110100101101001011010010110,
64'b1001011010010110100101101001011011110000111100001111000011110000,
64'b0011110011000011110000110011110000000000111111111111111100000000,
64'b0000111100001111111100001111000000110011110011000011001111001100,
64'b1100001100111100110000110011110010010110100101101001011010010110,
64'b0110100110010110011010011001011001011010101001011010010101011010,
64'b0011001111001100001100111100110011001100110011001100110011001100,
64'b0101101001011010010110100101101010100101101001010101101001011010,
64'b0110011001100110011001100110011000111100001111000011110000111100,
64'b1010010110100101010110100101101001100110100110011001100101100110,
64'b1111111100000000111111110000000011001100110011001100110011001100,
64'b1001011001101001011010011001011000000000111111111111111100000000,
64'b0110011010011001100110010110011001101001100101100110100110010110,
64'b1001100110011001011001100110011001101001100101100110100110010110,
64'b1100001100111100110000110011110011111111000000001111111100000000,
64'b1111000000001111000011111111000011111111111111110000000000000000,
64'b0101010110101010010101011010101010100101101001010101101001011010,
64'b0101101010100101101001010101101011000011001111001100001100111100,
64'b0011110011000011110000110011110011001100001100110011001111001100,
64'b1111000011110000111100001111000001011010010110100101101001011010,
64'b1001100101100110100110010110011000110011110011000011001111001100,
64'b0011110000111100001111000011110010100101010110101010010101011010,
64'b0011001111001100001100111100110011000011110000110011110000111100,
64'b0101010101010101101010101010101001011010010110100101101001011010,
64'b0011110011000011110000110011110011111111111111110000000000000000,
64'b0110100101101001100101101001011010010110011010010110100110010110,
64'b1001011010010110100101101001011000111100110000111100001100111100,
64'b0101101010100101101001010101101011111111111111110000000000000000,
64'b0000000011111111111111110000000000000000000000000000000000000000,
64'b1001100110011001011001100110011010011001011001101001100101100110,
64'b1100110000110011001100111100110001011010101001011010010101011010,
64'b0101101010100101101001010101101000001111000011111111000011110000,
64'b0101010110101010010101011010101010011001011001101001100101100110,
64'b1010101001010101010101011010101000001111111100000000111111110000,
64'b1100110011001100110011001100110001100110011001100110011001100110,
64'b1100110011001100110011001100110010100101010110101010010101011010,
64'b1001011001101001011010011001011011111111111111110000000000000000,
64'b1001100101100110100110010110011011000011110000110011110000111100,
64'b1010010101011010101001010101101001010101010101011010101010101010,
64'b1111000011110000111100001111000000001111111100000000111111110000,
64'b1100001100111100110000110011110001100110011001100110011001100110,
64'b1010101001010101010101011010101010010110100101101001011010010110,
64'b0011001100110011110011001100110001100110011001100110011001100110,
64'b1100001111000011001111000011110000000000000000000000000000000000,
64'b0000000011111111111111110000000011110000000011110000111111110000,
64'b0011001111001100001100111100110011111111000000001111111100000000,
64'b1001100101100110100110010110011000000000111111111111111100000000,
64'b1001011010010110100101101001011000111100001111000011110000111100,
64'b0011110000111100001111000011110011001100001100110011001111001100,
64'b1010101010101010101010101010101000000000000000000000000000000000,
64'b1111000000001111000011111111000010100101010110101010010101011010,
64'b0110100101101001100101101001011001100110011001100110011001100110,
64'b0000111111110000000011111111000010101010010101010101010110101010,
64'b0011001100110011110011001100110000111100001111000011110000111100,
64'b1001100101100110100110010110011011000011001111001100001100111100,
64'b0110100101101001100101101001011000111100001111000011110000111100,
64'b0110011010011001100110010110011000000000000000000000000000000000,
64'b0101010110101010010101011010101000000000111111111111111100000000,
64'b0110100110010110011010011001011010101010101010101010101010101010,
64'b1100001100111100110000110011110001010101010101011010101010101010,
64'b0000111111110000000011111111000010100101010110101010010101011010,
64'b1100001100111100110000110011110000001111000011111111000011110000,
64'b0101101010100101101001010101101010101010101010101010101010101010,
64'b1001100110011001011001100110011011001100001100110011001111001100,
64'b1100110011001100110011001100110000111100001111000011110000111100,
64'b0101101010100101101001010101101000110011001100111100110011001100,
64'b0011001111001100001100111100110010100101010110101010010101011010,
64'b1100001100111100110000110011110011110000000011110000111111110000,
64'b1111000000001111000011111111000000001111111100000000111111110000,
64'b1010101010101010101010101010101000000000000000000000000000000000,
64'b1001100101100110100110010110011011111111111111110000000000000000,
64'b1111000011110000111100001111000001100110011001100110011001100110,
64'b1111000000001111000011111111000011001100110011001100110011001100,
64'b0000000011111111111111110000000001100110100110011001100101100110,
64'b1111000000001111000011111111000011111111000000001111111100000000,
64'b1100110000110011001100111100110001100110011001100110011001100110,
64'b1001011010010110100101101001011000001111000011111111000011110000,
64'b0101101001011010010110100101101010100101010110101010010101011010,
64'b1100110000110011001100111100110011110000111100001111000011110000,
64'b1010010110100101010110100101101001100110100110011001100101100110,
64'b1111000000001111000011111111000000000000111111111111111100000000,
64'b0000000011111111111111110000000010101010010101010101010110101010,
64'b0110011001100110011001100110011000000000000000000000000000000000,
64'b1100001111000011001111000011110000000000000000000000000000000000,
64'b1111111100000000111111110000000010010110100101101001011010010110,
64'b0000000000000000000000000000000011110000111100001111000011110000,
64'b1001100110011001011001100110011011000011110000110011110000111100,
64'b0110011010011001100110010110011001010101010101011010101010101010,
64'b0011001111001100001100111100110000111100001111000011110000111100,
64'b1111000011110000111100001111000011111111000000001111111100000000,
64'b1001011010010110100101101001011001100110100110011001100101100110,
64'b1111111111111111000000000000000011111111000000001111111100000000,
64'b0101101001011010010110100101101011000011110000110011110000111100,
64'b0000000000000000000000000000000001010101010101011010101010101010,
64'b0110011001100110011001100110011010011001100110010110011001100110,
64'b0101010101010101101010101010101010101010101010101010101010101010,
64'b0000111100001111111100001111000000000000000000000000000000000000,
64'b1001100101100110100110010110011011000011001111001100001100111100,
64'b1010101001010101010101011010101001010101101010100101010110101010,
64'b1111000011110000111100001111000000001111111100000000111111110000,
64'b1010010110100101010110100101101001100110011001100110011001100110,
64'b0011001111001100001100111100110010100101010110101010010101011010,
64'b0110011001100110011001100110011011111111111111110000000000000000,
64'b0110011001100110011001100110011011000011110000110011110000111100,
64'b1111000011110000111100001111000001010101010101011010101010101010,
64'b0101101001011010010110100101101000001111111100000000111111110000,
64'b1010101001010101010101011010101001100110011001100110011001100110,
64'b0000111100001111111100001111000010010110100101101001011010010110,
64'b0000111100001111111100001111000001100110011001100110011001100110,
64'b0101010101010101101010101010101000000000000000000000000000000000,
64'b1010010101011010101001010101101000001111111100000000111111110000,
64'b1001100110011001011001100110011010011001011001101001100101100110,
64'b0101010110101010010101011010101011001100001100110011001111001100,
64'b0011001111001100001100111100110011110000111100001111000011110000,
64'b1010010110100101010110100101101001011010010110100101101001011010,
64'b0011110000111100001111000011110010011001011001101001100101100110,
64'b0011110000111100001111000011110000000000000000000000000000000000,
64'b1111111100000000111111110000000010010110100101101001011010010110,
64'b0011001111001100001100111100110001101001011010011001011010010110,
64'b0011001100110011110011001100110010010110011010010110100110010110,
64'b0101010110101010010101011010101011110000000011110000111111110000,
64'b0101010110101010010101011010101011111111111111110000000000000000,
64'b0110011001100110011001100110011000000000111111111111111100000000,
64'b1001100101100110100110010110011011001100110011001100110011001100,
64'b0011110011000011110000110011110001101001100101100110100110010110,
64'b0101010101010101101010101010101011000011110000110011110000111100,
64'b1100001111000011001111000011110010011001011001101001100101100110,
64'b1010010110100101010110100101101010100101101001010101101001011010,
64'b0011110000111100001111000011110001011010101001011010010101011010,
64'b1010101010101010101010101010101010100101010110101010010101011010,
64'b0000111100001111111100001111000000110011110011000011001111001100,
64'b1100110000110011001100111100110000000000000000000000000000000000,
64'b0101101010100101101001010101101000111100001111000011110000111100,
64'b1010101010101010101010101010101010011001011001101001100101100110,
64'b1111000011110000111100001111000001101001011010011001011010010110,
64'b0011110011000011110000110011110001010101101010100101010110101010,
64'b0000111111110000000011111111000001101001100101100110100110010110,
64'b1111000011110000111100001111000000111100110000111100001100111100,
64'b1010101010101010101010101010101000001111111100000000111111110000,
64'b0110100110010110011010011001011001101001011010011001011010010110,
64'b0000111100001111111100001111000000110011110011000011001111001100,
64'b0011110000111100001111000011110001100110100110011001100101100110,
64'b0110100110010110011010011001011001100110100110011001100101100110,
64'b0000111111110000000011111111000000001111000011111111000011110000,
64'b0110011010011001100110010110011000000000000000000000000000000000,
64'b1100110011001100110011001100110000001111111100000000111111110000,
64'b0101010101010101101010101010101011000011110000110011110000111100,
64'b0011110011000011110000110011110011000011001111001100001100111100,
64'b1111000011110000111100001111000010011001100110010110011001100110,
64'b0110011001100110011001100110011011000011001111001100001100111100,
64'b0101010110101010010101011010101011110000000011110000111111110000,
64'b1100110011001100110011001100110010101010010101010101010110101010,
64'b0011110011000011110000110011110011000011001111001100001100111100,
64'b1111111100000000111111110000000010100101101001010101101001011010,
64'b1010010101011010101001010101101011000011110000110011110000111100,
64'b0011110011000011110000110011110001101001011010011001011010010110,
64'b0000000011111111111111110000000001010101101010100101010110101010,
64'b1100001111000011001111000011110010101010101010101010101010101010,
64'b0101101001011010010110100101101000000000111111111111111100000000,
64'b1100110011001100110011001100110000001111111100000000111111110000,
64'b0101101010100101101001010101101001011010101001011010010101011010,
64'b0101010110101010010101011010101000111100001111000011110000111100,
64'b0011110000111100001111000011110010100101010110101010010101011010,
64'b0011001111001100001100111100110010101010101010101010101010101010,
64'b0011110000111100001111000011110001010101010101011010101010101010,
64'b0011110011000011110000110011110010010110011010010110100110010110,
64'b1100001100111100110000110011110010100101101001010101101001011010,
64'b0101010101010101101010101010101000111100001111000011110000111100,
64'b0101010101010101101010101010101011001100110011001100110011001100,
64'b1010010110100101010110100101101001101001011010011001011010010110,
64'b0110011001100110011001100110011000001111111100000000111111110000,
64'b0011001100110011110011001100110001010101101010100101010110101010,
64'b1100001111000011001111000011110010011001011001101001100101100110,
64'b0000111111110000000011111111000000001111111100000000111111110000,
64'b1001100101100110100110010110011010100101101001010101101001011010,
64'b0011110000111100001111000011110000000000000000000000000000000000,
64'b1010010101011010101001010101101011001100110011001100110011001100,
64'b1100001100111100110000110011110011001100110011001100110011001100,
64'b0011110011000011110000110011110010010110011010010110100110010110,
64'b1100110011001100110011001100110010011001011001101001100101100110,
64'b0101010110101010010101011010101010100101010110101010010101011010,
64'b1100001100111100110000110011110011110000111100001111000011110000,
64'b0110100110010110011010011001011011000011001111001100001100111100,
64'b0101010110101010010101011010101010101010010101010101010110101010,
64'b0101101010100101101001010101101000110011001100111100110011001100,
64'b1001011001101001011010011001011011000011110000110011110000111100,
64'b0110100110010110011010011001011000000000111111111111111100000000,
64'b1100001100111100110000110011110000110011110011000011001111001100,
64'b0011110000111100001111000011110010101010101010101010101010101010,
64'b0110011001100110011001100110011001011010010110100101101001011010,
64'b0011110011000011110000110011110011110000111100001111000011110000,
64'b0011110011000011110000110011110000111100110000111100001100111100,
64'b1100110000110011001100111100110001101001011010011001011010010110,
64'b1010101001010101010101011010101011001100001100110011001111001100,
64'b0101010101010101101010101010101011111111000000001111111100000000,
64'b1100110000110011001100111100110011110000000011110000111111110000,
64'b1111000000001111000011111111000000110011001100111100110011001100,
64'b0110011001100110011001100110011001011010010110100101101001011010,
64'b1010010101011010101001010101101010100101010110101010010101011010,
64'b0101010110101010010101011010101001010101010101011010101010101010,
64'b1111000011110000111100001111000010100101101001010101101001011010,
64'b0011110000111100001111000011110011001100110011001100110011001100,
64'b0011110000111100001111000011110010011001011001101001100101100110,
64'b1111000000001111000011111111000011111111000000001111111100000000,
64'b0101101010100101101001010101101011110000000011110000111111110000,
64'b1010010110100101010110100101101001101001100101100110100110010110,
64'b1001100110011001011001100110011010100101101001010101101001011010,
64'b0110011001100110011001100110011001010101010101011010101010101010,
64'b1010010110100101010110100101101000000000111111111111111100000000,
64'b1010101001010101010101011010101001011010010110100101101001011010,
64'b1001011010010110100101101001011010011001011001101001100101100110,
64'b1100110000110011001100111100110011001100001100110011001111001100,
64'b0011001100110011110011001100110011001100110011001100110011001100,
64'b1111111100000000111111110000000010011001011001101001100101100110,
64'b0000111111110000000011111111000001011010010110100101101001011010,
64'b1010010101011010101001010101101011000011110000110011110000111100,
64'b0000000011111111111111110000000011111111111111110000000000000000,
64'b0110011010011001100110010110011000000000111111111111111100000000,
64'b1001100101100110100110010110011010010110011010010110100110010110,
64'b1001011010010110100101101001011000110011110011000011001111001100,
64'b1001011010010110100101101001011001100110011001100110011001100110,
64'b0011001111001100001100111100110001010101010101011010101010101010,
64'b1001100110011001011001100110011010011001011001101001100101100110,
64'b0110100110010110011010011001011011000011110000110011110000111100,
64'b0000111100001111111100001111000000001111000011111111000011110000,
64'b0101101001011010010110100101101001011010010110100101101001011010,
64'b0101010101010101101010101010101011000011110000110011110000111100,
64'b1111111100000000111111110000000000110011110011000011001111001100,
64'b1100110000110011001100111100110000001111111100000000111111110000,
64'b1111111111111111000000000000000010101010101010101010101010101010,
64'b0110100101101001100101101001011001010101010101011010101010101010,
64'b0110100101101001100101101001011010010110011010010110100110010110,
64'b1100001100111100110000110011110010100101101001010101101001011010,
64'b1100001100111100110000110011110000111100001111000011110000111100,
64'b0000111100001111111100001111000011001100110011001100110011001100,
64'b0011110000111100001111000011110001101001011010011001011010010110,
64'b1001011001101001011010011001011000001111111100000000111111110000,
64'b1111111100000000111111110000000001010101101010100101010110101010,
64'b1001100101100110100110010110011010011001011001101001100101100110,
64'b1100110011001100110011001100110000001111111100000000111111110000,
64'b1010101010101010101010101010101001011010010110100101101001011010,
64'b1100110011001100110011001100110011110000111100001111000011110000,
64'b0011001111001100001100111100110001011010010110100101101001011010,
64'b0000111100001111111100001111000001011010010110100101101001011010,
64'b1100001100111100110000110011110001011010010110100101101001011010,
64'b0101010110101010010101011010101011111111111111110000000000000000,
64'b1010101010101010101010101010101001100110011001100110011001100110,
64'b1010010110100101010110100101101010011001011001101001100101100110,
64'b0110011010011001100110010110011011000011001111001100001100111100,
64'b1001011001101001011010011001011011110000111100001111000011110000,
64'b0110100110010110011010011001011001101001100101100110100110010110,
64'b0110011001100110011001100110011010100101101001010101101001011010,
64'b1100001111000011001111000011110010101010101010101010101010101010,
64'b0000000000000000000000000000000000001111111100000000111111110000,
64'b1001011010010110100101101001011001010101101010100101010110101010,
64'b0011110011000011110000110011110000110011110011000011001111001100,
64'b1111000000001111000011111111000000110011110011000011001111001100,
64'b1001100110011001011001100110011000110011110011000011001111001100,
64'b0110011010011001100110010110011000000000000000000000000000000000,
64'b0110011001100110011001100110011010010110100101101001011010010110,
64'b1001011001101001011010011001011011000011110000110011110000111100,
64'b0000111111110000000011111111000011110000000011110000111111110000,
64'b0000000000000000000000000000000011111111000000001111111100000000,
64'b1111111111111111000000000000000000111100110000111100001100111100,
64'b0101101001011010010110100101101000110011110011000011001111001100,
64'b1100110000110011001100111100110001100110011001100110011001100110,
64'b1010101010101010101010101010101011111111000000001111111100000000,
64'b1010010101011010101001010101101000110011001100111100110011001100,
64'b1100001111000011001111000011110000001111000011111111000011110000,
64'b1010010101011010101001010101101000001111000011111111000011110000,
64'b0101010110101010010101011010101000001111000011111111000011110000,
64'b0011110011000011110000110011110000000000000000000000000000000000,
64'b0011110000111100001111000011110011000011001111001100001100111100,
64'b1001100101100110100110010110011000001111111100000000111111110000,
64'b1100110011001100110011001100110010101010010101010101010110101010,
64'b1001011001101001011010011001011001010101010101011010101010101010,
64'b0110100110010110011010011001011011110000000011110000111111110000,
64'b1111111100000000111111110000000010100101101001010101101001011010,
64'b1100110011001100110011001100110000111100001111000011110000111100,
64'b0110011001100110011001100110011000000000000000000000000000000000,
64'b1100110000110011001100111100110011110000111100001111000011110000,
64'b0000111111110000000011111111000001010101101010100101010110101010,
64'b0110011010011001100110010110011001010101101010100101010110101010,
64'b0011001100110011110011001100110001010101101010100101010110101010,
64'b1111000000001111000011111111000010101010101010101010101010101010,
64'b1010010101011010101001010101101011110000000011110000111111110000,
64'b1100001111000011001111000011110000000000111111111111111100000000,
64'b1111000011110000111100001111000000110011001100111100110011001100,
64'b0011110011000011110000110011110001100110011001100110011001100110,
64'b1001011001101001011010011001011010101010010101010101010110101010,
64'b1111111111111111000000000000000010011001011001101001100101100110,
64'b1111000011110000111100001111000010100101010110101010010101011010,
64'b0011110000111100001111000011110000000000000000000000000000000000,
64'b0110100101101001100101101001011011111111000000001111111100000000,
64'b1001100110011001011001100110011000110011001100111100110011001100,
64'b1100110011001100110011001100110000110011001100111100110011001100,
64'b1001100101100110100110010110011000110011001100111100110011001100,
64'b1111111111111111000000000000000011001100110011001100110011001100,
64'b1100110000110011001100111100110000000000111111111111111100000000,
64'b1010101001010101010101011010101001010101010101011010101010101010,
64'b0011001100110011110011001100110001011010010110100101101001011010,
64'b0110011001100110011001100110011010010110100101101001011010010110,
64'b1111111111111111000000000000000000110011001100111100110011001100,
64'b1100110011001100110011001100110001101001011010011001011010010110,
64'b1001011001101001011010011001011011001100001100110011001111001100,
64'b0000111111110000000011111111000000000000000000000000000000000000,
64'b1010010101011010101001010101101001010101010101011010101010101010,
64'b1010010101011010101001010101101011110000111100001111000011110000,
64'b0101010101010101101010101010101001011010010110100101101001011010,
64'b0000000011111111111111110000000001011010010110100101101001011010,
64'b0101010110101010010101011010101001011010010110100101101001011010,
64'b0000111100001111111100001111000011111111111111110000000000000000,
64'b0011110000111100001111000011110001100110011001100110011001100110,
64'b0011110011000011110000110011110010011001011001101001100101100110,
64'b0000000011111111111111110000000011000011001111001100001100111100,
64'b0110100110010110011010011001011011110000111100001111000011110000,
64'b0011110000111100001111000011110001101001100101100110100110010110,
64'b1111111100000000111111110000000010100101101001010101101001011010,
64'b0101010110101010010101011010101010101010101010101010101010101010,
64'b0110011010011001100110010110011010101010101010101010101010101010,
64'b1100110000110011001100111100110001100110011001100110011001100110,
64'b1100110011001100110011001100110000111100110000111100001100111100,
64'b0101010101010101101010101010101011110000111100001111000011110000,
64'b1001100110011001011001100110011001100110011001100110011001100110,
64'b1111111100000000111111110000000010101010101010101010101010101010,
64'b1010010101011010101001010101101000110011001100111100110011001100,
64'b1111000000001111000011111111000010100101010110101010010101011010,
64'b0101010101010101101010101010101001100110011001100110011001100110,
64'b1001011001101001011010011001011010010110100101101001011010010110,
64'b0000111111110000000011111111000001011010101001011010010101011010,
64'b1111111111111111000000000000000011110000000011110000111111110000,
64'b1100110011001100110011001100110001100110011001100110011001100110,
64'b1010010110100101010110100101101000000000000000000000000000000000,
64'b1001011001101001011010011001011000001111111100000000111111110000,
64'b0101010101010101101010101010101011111111000000001111111100000000,
64'b0000111111110000000011111111000010010110100101101001011010010110,
64'b1100001100111100110000110011110001101001100101100110100110010110,
64'b1111111111111111000000000000000001100110011001100110011001100110,
64'b0110100110010110011010011001011001010101010101011010101010101010,
64'b0110011001100110011001100110011000000000000000000000000000000000,
64'b1111000000001111000011111111000010101010010101010101010110101010,
64'b1111111111111111000000000000000010101010101010101010101010101010,
64'b1100110000110011001100111100110010101010010101010101010110101010,
64'b1100001111000011001111000011110001101001100101100110100110010110,
64'b0101101001011010010110100101101010010110100101101001011010010110,
64'b0101010110101010010101011010101010101010101010101010101010101010,
64'b1010010110100101010110100101101000000000111111111111111100000000,
64'b0110100101101001100101101001011011111111111111110000000000000000,
64'b0110100101101001100101101001011011000011001111001100001100111100,
64'b1010010110100101010110100101101000111100110000111100001100111100,
64'b1010101010101010101010101010101000111100001111000011110000111100,
64'b0011001111001100001100111100110011001100110011001100110011001100,
64'b0101101010100101101001010101101010101010101010101010101010101010,
64'b1001011010010110100101101001011000110011001100111100110011001100,
64'b1100001100111100110000110011110001100110011001100110011001100110,
64'b1100001111000011001111000011110000110011001100111100110011001100,
64'b0110011010011001100110010110011010010110011010010110100110010110,
64'b1001100101100110100110010110011011000011001111001100001100111100,
64'b0011001100110011110011001100110001100110011001100110011001100110,
64'b0011001111001100001100111100110011111111111111110000000000000000,
64'b0110100110010110011010011001011010101010101010101010101010101010,
64'b0110100110010110011010011001011001011010101001011010010101011010,
64'b1001100101100110100110010110011011110000000011110000111111110000,
64'b0110011001100110011001100110011010100101010110101010010101011010,
64'b0000111100001111111100001111000011110000111100001111000011110000,
64'b1100110000110011001100111100110011001100110011001100110011001100,
64'b0110100110010110011010011001011011110000111100001111000011110000,
64'b1111000000001111000011111111000010010110100101101001011010010110,
64'b0000111111110000000011111111000011110000111100001111000011110000,
64'b0110100101101001100101101001011010010110011010010110100110010110,
64'b1001011010010110100101101001011010100101010110101010010101011010,
64'b0011110000111100001111000011110001011010010110100101101001011010,
64'b1001011001101001011010011001011000110011110011000011001111001100,
64'b0011001111001100001100111100110001101001011010011001011010010110,
64'b1111111111111111000000000000000000001111000011111111000011110000,
64'b1001011001101001011010011001011011111111111111110000000000000000,
64'b1001011010010110100101101001011011001100001100110011001111001100,
64'b0101101010100101101001010101101001011010101001011010010101011010,
64'b1100001100111100110000110011110010010110011010010110100110010110,
64'b0000000000000000000000000000000001101001011010011001011010010110,
64'b0110100101101001100101101001011010101010101010101010101010101010,
64'b1100110000110011001100111100110010011001011001101001100101100110,
64'b0000000011111111111111110000000011111111000000001111111100000000,
64'b0110100110010110011010011001011010011001011001101001100101100110,
64'b1100001100111100110000110011110000110011110011000011001111001100,
64'b0000111100001111111100001111000000001111000011111111000011110000,
64'b1010101010101010101010101010101011000011001111001100001100111100,
64'b1100001100111100110000110011110001010101101010100101010110101010,
64'b1100001111000011001111000011110010101010101010101010101010101010,
64'b1100001100111100110000110011110010100101101001010101101001011010,
64'b0110100110010110011010011001011001100110100110011001100101100110,
64'b0011110000111100001111000011110010010110011010010110100110010110,
64'b1001011001101001011010011001011001101001100101100110100110010110,
64'b1010101010101010101010101010101001100110011001100110011001100110,
64'b1100001111000011001111000011110011000011110000110011110000111100,
64'b1001011010010110100101101001011011111111111111110000000000000000,
64'b0110100110010110011010011001011000111100001111000011110000111100,
64'b0011110011000011110000110011110000001111000011111111000011110000,
64'b1100110011001100110011001100110011111111000000001111111100000000,
64'b0110100101101001100101101001011001011010101001011010010101011010,
64'b0011001100110011110011001100110000110011001100111100110011001100,
64'b0101101001011010010110100101101011001100110011001100110011001100,
64'b1111000000001111000011111111000000110011110011000011001111001100,
64'b1001100101100110100110010110011001101001011010011001011010010110,
64'b0110100101101001100101101001011010010110011010010110100110010110,
64'b1010101010101010101010101010101010010110011010010110100110010110,
64'b0000111111110000000011111111000000111100001111000011110000111100,
64'b0110100110010110011010011001011000001111111100000000111111110000,
64'b1010101001010101010101011010101010101010101010101010101010101010,
64'b1100001100111100110000110011110010100101010110101010010101011010,
64'b1111000000001111000011111111000011111111000000001111111100000000,
64'b0101101001011010010110100101101001010101010101011010101010101010,
64'b1100001100111100110000110011110011001100001100110011001111001100,
64'b0101101001011010010110100101101001011010010110100101101001011010,
64'b1001100101100110100110010110011001011010010110100101101001011010,
64'b0000000011111111111111110000000000001111000011111111000011110000,
64'b0110100101101001100101101001011011000011001111001100001100111100,
64'b1100001100111100110000110011110010010110011010010110100110010110,
64'b0110011001100110011001100110011010010110011010010110100110010110,
64'b0000000011111111111111110000000010100101010110101010010101011010,
64'b0011110011000011110000110011110000000000111111111111111100000000,
64'b0011001100110011110011001100110011001100110011001100110011001100,
64'b1010010101011010101001010101101000110011110011000011001111001100,
64'b1010101001010101010101011010101011111111111111110000000000000000,
64'b1001100101100110100110010110011011001100110011001100110011001100,
64'b1111000000001111000011111111000010100101101001010101101001011010,
64'b0011001111001100001100111100110010011001011001101001100101100110,
64'b1100001111000011001111000011110000110011110011000011001111001100,
64'b1111111111111111000000000000000011111111000000001111111100000000,
64'b0110100110010110011010011001011001011010101001011010010101011010,
64'b0101101010100101101001010101101000111100110000111100001100111100,
64'b0011110000111100001111000011110010010110011010010110100110010110,
64'b1111111111111111000000000000000001100110100110011001100101100110,
64'b0101101010100101101001010101101011111111111111110000000000000000,
64'b0101101001011010010110100101101001011010010110100101101001011010,
64'b1001100101100110100110010110011011110000111100001111000011110000,
64'b1001100110011001011001100110011010101010101010101010101010101010,
64'b0110100101101001100101101001011001011010010110100101101001011010,
64'b0000000011111111111111110000000000110011110011000011001111001100,
64'b1010010110100101010110100101101001101001011010011001011010010110,
64'b0000111111110000000011111111000000001111000011111111000011110000,
64'b1010101010101010101010101010101011111111111111110000000000000000,
64'b1001011001101001011010011001011011001100001100110011001111001100,
64'b1100110000110011001100111100110001011010101001011010010101011010,
64'b1010010101011010101001010101101010010110011010010110100110010110,
64'b0000000000000000000000000000000001101001011010011001011010010110,
64'b0110011010011001100110010110011010101010101010101010101010101010,
64'b1001100101100110100110010110011010011001011001101001100101100110,
64'b0011110000111100001111000011110011111111000000001111111100000000,
64'b1010010101011010101001010101101001100110011001100110011001100110,
64'b1010010101011010101001010101101001010101010101011010101010101010,
64'b0101010101010101101010101010101011111111111111110000000000000000,
64'b0011110011000011110000110011110011000011110000110011110000111100,
64'b0011110000111100001111000011110011111111111111110000000000000000,
64'b0101101010100101101001010101101010101010101010101010101010101010,
64'b1100110011001100110011001100110010011001011001101001100101100110,
64'b0110100101101001100101101001011011000011001111001100001100111100,
64'b0011110011000011110000110011110011001100110011001100110011001100,
64'b0110100101101001100101101001011001010101010101011010101010101010,
64'b0011001100110011110011001100110000001111000011111111000011110000,
64'b0101101010100101101001010101101010101010101010101010101010101010,
64'b1100110011001100110011001100110001100110011001100110011001100110,
64'b0110100101101001100101101001011010010110100101101001011010010110,
64'b0110100101101001100101101001011011001100110011001100110011001100,
64'b1001100110011001011001100110011010101010101010101010101010101010,
64'b0110011001100110011001100110011010100101010110101010010101011010,
64'b1001100101100110100110010110011010101010101010101010101010101010,
64'b1001011010010110100101101001011001100110011001100110011001100110,
64'b1001011010010110100101101001011011000011110000110011110000111100,
64'b1010101001010101010101011010101011110000000011110000111111110000,
64'b0110011001100110011001100110011011110000111100001111000011110000,
64'b0000000011111111111111110000000011001100110011001100110011001100,
64'b0110100101101001100101101001011001010101101010100101010110101010,
64'b0011110000111100001111000011110001100110011001100110011001100110,
64'b1001011010010110100101101001011000111100001111000011110000111100,
64'b0110011001100110011001100110011001101001100101100110100110010110,
64'b1100110011001100110011001100110011110000111100001111000011110000,
64'b1100001111000011001111000011110011001100110011001100110011001100,
64'b1010101001010101010101011010101011001100001100110011001111001100,
64'b1111111111111111000000000000000011001100110011001100110011001100,
64'b1001100110011001011001100110011000111100001111000011110000111100,
64'b0000111111110000000011111111000000001111111100000000111111110000,
64'b0101101001011010010110100101101010101010010101010101010110101010,
64'b1010101001010101010101011010101001010101101010100101010110101010,
64'b1001011010010110100101101001011011110000111100001111000011110000,
64'b0101101010100101101001010101101000110011001100111100110011001100,
64'b1111111111111111000000000000000000111100001111000011110000111100,
64'b0000111111110000000011111111000000001111111100000000111111110000,
64'b0011110000111100001111000011110000111100110000111100001100111100,
64'b1111000011110000111100001111000011111111000000001111111100000000,
64'b0000111111110000000011111111000011110000111100001111000011110000,
64'b1001100110011001011001100110011000001111000011111111000011110000,
64'b1010101010101010101010101010101001011010010110100101101001011010,
64'b1001011010010110100101101001011000001111111100000000111111110000,
64'b1010101001010101010101011010101000000000111111111111111100000000,
64'b0011001111001100001100111100110000110011001100111100110011001100,
64'b0011001100110011110011001100110010011001100110010110011001100110,
64'b0110100110010110011010011001011011111111000000001111111100000000,
64'b1100110000110011001100111100110011110000111100001111000011110000,
64'b1010101010101010101010101010101010100101010110101010010101011010,
64'b0101010110101010010101011010101011111111000000001111111100000000,
64'b1010101010101010101010101010101011110000000011110000111111110000,
64'b0101101001011010010110100101101001010101010101011010101010101010,
64'b0101010110101010010101011010101011111111000000001111111100000000,
64'b0000000011111111111111110000000011111111000000001111111100000000,
64'b0101101001011010010110100101101010011001011001101001100101100110,
64'b1001100110011001011001100110011000000000111111111111111100000000,
64'b1111111111111111000000000000000011111111111111110000000000000000,
64'b1100110011001100110011001100110001011010010110100101101001011010,
64'b1100110000110011001100111100110010010110100101101001011010010110,
64'b1111111100000000111111110000000001010101010101011010101010101010,
64'b0011110000111100001111000011110011111111000000001111111100000000,
64'b0011110011000011110000110011110011001100001100110011001111001100,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1100001100111100110000110011110000000000111111111111111100000000,
64'b1001011010010110100101101001011001100110011001100110011001100110,
64'b0110011001100110011001100110011001010101010101011010101010101010,
64'b1100001100111100110000110011110011111111111111110000000000000000,
64'b1010010101011010101001010101101011000011110000110011110000111100,
64'b0110011010011001100110010110011011111111111111110000000000000000,
64'b0110011001100110011001100110011010101010101010101010101010101010,
64'b0011001100110011110011001100110010011001011001101001100101100110,
64'b0011001111001100001100111100110011000011001111001100001100111100,
64'b0011110000111100001111000011110011001100110011001100110011001100,
64'b0011110011000011110000110011110001010101010101011010101010101010,
64'b1010101010101010101010101010101000001111000011111111000011110000,
64'b0110011001100110011001100110011010101010101010101010101010101010,
64'b0101101010100101101001010101101001011010101001011010010101011010,
64'b1100001100111100110000110011110000110011110011000011001111001100,
64'b0011110000111100001111000011110010011001100110010110011001100110,
64'b1111000000001111000011111111000010010110011010010110100110010110,
64'b1100110000110011001100111100110010011001011001101001100101100110,
64'b1100001111000011001111000011110011110000000011110000111111110000,
64'b1001011010010110100101101001011010101010101010101010101010101010,
64'b1111000011110000111100001111000010101010101010101010101010101010,
64'b1010010110100101010110100101101011001100110011001100110011001100,
64'b0000111111110000000011111111000010011001100110010110011001100110,
64'b1111000000001111000011111111000011111111111111110000000000000000,
64'b0110011001100110011001100110011000001111000011111111000011110000,
64'b0011110000111100001111000011110010101010101010101010101010101010,
64'b0110100101101001100101101001011001101001011010011001011010010110,
64'b1111111111111111000000000000000000000000111111111111111100000000,
64'b0101101010100101101001010101101001101001011010011001011010010110,
64'b0011110000111100001111000011110010101010101010101010101010101010,
64'b1001100110011001011001100110011001010101010101011010101010101010,
64'b1111111111111111000000000000000001011010010110100101101001011010,
64'b1010010101011010101001010101101010101010101010101010101010101010,
64'b1001011001101001011010011001011010100101101001010101101001011010,
64'b0000111100001111111100001111000011001100001100110011001111001100,
64'b1100001100111100110000110011110001010101010101011010101010101010,
64'b0011001111001100001100111100110010011001100110010110011001100110,
64'b1100110000110011001100111100110000001111000011111111000011110000,
64'b1100001100111100110000110011110010101010101010101010101010101010,
64'b0110011001100110011001100110011011000011001111001100001100111100,
64'b0000111111110000000011111111000001010101010101011010101010101010,
64'b0011001111001100001100111100110001101001100101100110100110010110,
64'b1001100110011001011001100110011001100110011001100110011001100110,
64'b0000000000000000000000000000000011001100110011001100110011001100,
64'b1111000000001111000011111111000010011001011001101001100101100110,
64'b1010101001010101010101011010101011001100110011001100110011001100,
64'b0101010110101010010101011010101000110011110011000011001111001100,
64'b0110100101101001100101101001011010100101101001010101101001011010,
64'b0011001111001100001100111100110001100110011001100110011001100110,
64'b0011110000111100001111000011110010010110100101101001011010010110,
64'b0101010110101010010101011010101001010101101010100101010110101010,
64'b0110100110010110011010011001011001100110011001100110011001100110,
64'b1001011010010110100101101001011001011010101001011010010101011010,
64'b0000000011111111111111110000000011001100110011001100110011001100,
64'b0000111100001111111100001111000010010110011010010110100110010110,
64'b0011110000111100001111000011110000111100001111000011110000111100,
64'b1010101010101010101010101010101011110000111100001111000011110000,
64'b0000000011111111111111110000000011000011110000110011110000111100,
64'b1001100110011001011001100110011011110000111100001111000011110000,
64'b1001100110011001011001100110011000001111000011111111000011110000,
64'b1100001100111100110000110011110000110011110011000011001111001100,
64'b1010010110100101010110100101101010010110100101101001011010010110,
64'b0000111111110000000011111111000011000011001111001100001100111100,
64'b0011001100110011110011001100110000110011001100111100110011001100,
64'b1100001100111100110000110011110000111100001111000011110000111100,
64'b0110011001100110011001100110011011000011110000110011110000111100,
64'b0101101010100101101001010101101011111111000000001111111100000000,
64'b0000000011111111111111110000000001101001100101100110100110010110,
64'b1001100110011001011001100110011010011001100110010110011001100110,
64'b1111000011110000111100001111000011000011001111001100001100111100,
64'b1010010101011010101001010101101001010101010101011010101010101010,
64'b0101101001011010010110100101101010011001011001101001100101100110,
64'b1111111111111111000000000000000010010110011010010110100110010110,
64'b0110011001100110011001100110011010011001011001101001100101100110,
64'b0101101010100101101001010101101010101010010101010101010110101010,
64'b1001100101100110100110010110011011000011001111001100001100111100,
64'b1010101001010101010101011010101010101010010101010101010110101010,
64'b0110100110010110011010011001011001101001100101100110100110010110,
64'b0011001111001100001100111100110010100101010110101010010101011010,
64'b0110100101101001100101101001011001010101010101011010101010101010,
64'b0000000000000000000000000000000000111100110000111100001100111100,
64'b1010101001010101010101011010101000111100001111000011110000111100,
64'b0110100110010110011010011001011001011010101001011010010101011010,
64'b1001011010010110100101101001011011001100110011001100110011001100,
64'b1111111100000000111111110000000001101001011010011001011010010110,
64'b0110100101101001100101101001011000111100110000111100001100111100,
64'b1010101001010101010101011010101001101001011010011001011010010110,
64'b1010010101011010101001010101101000110011001100111100110011001100,
64'b0101101001011010010110100101101001011010101001011010010101011010,
64'b0110100110010110011010011001011000110011001100111100110011001100,
64'b1010010101011010101001010101101001101001100101100110100110010110,
64'b0000000011111111111111110000000011001100001100110011001111001100,
64'b0110011001100110011001100110011011001100110011001100110011001100,
64'b1111111111111111000000000000000001011010101001011010010101011010,
64'b0000111111110000000011111111000010100101010110101010010101011010,
64'b1010101001010101010101011010101011001100001100110011001111001100,
64'b1001100110011001011001100110011001011010010110100101101001011010,
64'b0011001100110011110011001100110011000011001111001100001100111100,
64'b1010101001010101010101011010101001011010101001011010010101011010,
64'b1010010101011010101001010101101001101001100101100110100110010110,
64'b0000111111110000000011111111000001011010010110100101101001011010,
64'b0000000011111111111111110000000001100110100110011001100101100110,
64'b0110011001100110011001100110011001011010010110100101101001011010,
64'b1111111100000000111111110000000001101001100101100110100110010110,
64'b0101010101010101101010101010101010100101101001010101101001011010,
64'b1001011010010110100101101001011001011010010110100101101001011010,
64'b0000000000000000000000000000000011001100001100110011001111001100,
64'b1010101001010101010101011010101001100110100110011001100101100110,
64'b0011001100110011110011001100110000001111000011111111000011110000,
64'b1001011010010110100101101001011010011001011001101001100101100110,
64'b0101101001011010010110100101101011110000000011110000111111110000,
64'b1001100110011001011001100110011011001100001100110011001111001100,
64'b0110011010011001100110010110011010010110011010010110100110010110,
64'b0000000011111111111111110000000000110011110011000011001111001100,
64'b1111111111111111000000000000000011000011110000110011110000111100,
64'b1001011010010110100101101001011010011001011001101001100101100110,
64'b0000000000000000000000000000000011000011001111001100001100111100,
64'b0110011001100110011001100110011010011001011001101001100101100110,
64'b0110100110010110011010011001011010011001011001101001100101100110,
64'b0000000000000000000000000000000000001111000011111111000011110000,
64'b0011001100110011110011001100110001101001011010011001011010010110,
64'b0101101001011010010110100101101001010101101010100101010110101010,
64'b0110100110010110011010011001011001101001011010011001011010010110,
64'b0011001111001100001100111100110000000000111111111111111100000000,
64'b0011110000111100001111000011110010100101101001010101101001011010,
64'b0110100101101001100101101001011010010110011010010110100110010110,
64'b0101010101010101101010101010101010100101101001010101101001011010,
64'b1010101010101010101010101010101000001111111100000000111111110000,
64'b0110100110010110011010011001011001101001011010011001011010010110,
64'b0000000000000000000000000000000000001111111100000000111111110000,
64'b1001011010010110100101101001011011000011110000110011110000111100,
64'b0011110011000011110000110011110011000011110000110011110000111100,
64'b0000000000000000000000000000000011111111000000001111111100000000,
64'b1111000011110000111100001111000001101001100101100110100110010110,
64'b1001100101100110100110010110011010011001100110010110011001100110,
64'b0011110011000011110000110011110011000011001111001100001100111100,
64'b0000111100001111111100001111000001010101010101011010101010101010,
64'b0000111111110000000011111111000010011001011001101001100101100110,
64'b1100001100111100110000110011110010010110011010010110100110010110,
64'b0110011001100110011001100110011010011001011001101001100101100110,
64'b0110011001100110011001100110011010101010010101010101010110101010,
64'b0011110011000011110000110011110011000011001111001100001100111100,
64'b0000000000000000000000000000000001010101101010100101010110101010,
64'b1001011001101001011010011001011001101001011010011001011010010110,
64'b0110100110010110011010011001011011000011110000110011110000111100,
64'b1001100110011001011001100110011000110011110011000011001111001100,
64'b1111111111111111000000000000000000111100110000111100001100111100,
64'b1100001111000011001111000011110011000011001111001100001100111100,
64'b0000000000000000000000000000000010011001100110010110011001100110,
64'b0000000000000000000000000000000010101010101010101010101010101010,
64'b0101101010100101101001010101101000111100110000111100001100111100,
64'b0000111111110000000011111111000011110000000011110000111111110000,
64'b0101010110101010010101011010101001011010101001011010010101011010,
64'b0000111100001111111100001111000010100101101001010101101001011010,
64'b1111000000001111000011111111000000000000111111111111111100000000,
64'b0000111111110000000011111111000011000011001111001100001100111100,
64'b1010101010101010101010101010101011000011001111001100001100111100,
64'b1111111111111111000000000000000010100101010110101010010101011010,
64'b1010010110100101010110100101101010100101101001010101101001011010,
64'b0101010101010101101010101010101011110000000011110000111111110000,
64'b0110011010011001100110010110011001011010101001011010010101011010,
64'b1010101010101010101010101010101000111100001111000011110000111100,
64'b0000000000000000000000000000000001100110011001100110011001100110,
64'b1001011010010110100101101001011011110000000011110000111111110000,
64'b1010010110100101010110100101101010101010010101010101010110101010,
64'b0110011010011001100110010110011001100110100110011001100101100110,
64'b1111000000001111000011111111000010011001011001101001100101100110,
64'b0101101001011010010110100101101001010101010101011010101010101010,
64'b0101101001011010010110100101101010100101010110101010010101011010,
64'b0101101010100101101001010101101011110000000011110000111111110000,
64'b0110100110010110011010011001011011001100001100110011001111001100,
64'b0000000011111111111111110000000000110011110011000011001111001100,
64'b1001100110011001011001100110011010101010010101010101010110101010,
64'b1010101010101010101010101010101001100110100110011001100101100110,
64'b0110011001100110011001100110011010100101010110101010010101011010,
64'b0000000000000000000000000000000000111100001111000011110000111100,
64'b1001100110011001011001100110011000000000111111111111111100000000,
64'b0011110000111100001111000011110010011001100110010110011001100110,
64'b0011110011000011110000110011110001101001011010011001011010010110,
64'b1010010101011010101001010101101001101001011010011001011010010110,
64'b0110100101101001100101101001011011001100110011001100110011001100,
64'b0011110000111100001111000011110010011001011001101001100101100110,
64'b0110011010011001100110010110011010101010010101010101010110101010,
64'b1001011001101001011010011001011010100101101001010101101001011010,
64'b1111111111111111000000000000000010100101101001010101101001011010,
64'b1001011010010110100101101001011000110011001100111100110011001100,
64'b0110011001100110011001100110011001101001011010011001011010010110,
64'b0011110000111100001111000011110001100110100110011001100101100110,
64'b0000000000000000000000000000000000001111111100000000111111110000,
64'b0011110000111100001111000011110011111111111111110000000000000000,
64'b1010010101011010101001010101101010010110100101101001011010010110,
64'b1111000000001111000011111111000001101001100101100110100110010110,
64'b0110011010011001100110010110011001101001100101100110100110010110,
64'b1100001100111100110000110011110001011010010110100101101001011010,
64'b1010010101011010101001010101101000111100001111000011110000111100,
64'b1111111100000000111111110000000010011001100110010110011001100110,
64'b1111111111111111000000000000000010011001011001101001100101100110,
64'b0011001100110011110011001100110010011001011001101001100101100110,
64'b1001011001101001011010011001011001011010010110100101101001011010,
64'b1111111111111111000000000000000001101001100101100110100110010110,
64'b0000111111110000000011111111000001101001011010011001011010010110,
64'b0000000000000000000000000000000010101010010101010101010110101010,
64'b0101010101010101101010101010101000000000000000000000000000000000,
64'b1100001111000011001111000011110001101001100101100110100110010110,
64'b0101010101010101101010101010101000111100110000111100001100111100,
64'b0110011001100110011001100110011000111100110000111100001100111100,
64'b1010101010101010101010101010101000110011110011000011001111001100,
64'b0011110000111100001111000011110000001111111100000000111111110000,
64'b0110100110010110011010011001011000111100001111000011110000111100,
64'b0110100110010110011010011001011001101001011010011001011010010110,
64'b1100001111000011001111000011110011000011110000110011110000111100,
64'b0110100110010110011010011001011000110011110011000011001111001100,
64'b0110100101101001100101101001011000111100110000111100001100111100,
64'b1010101001010101010101011010101011000011001111001100001100111100,
64'b0000000000000000000000000000000010011001100110010110011001100110,
64'b1001011001101001011010011001011010101010101010101010101010101010,
64'b1010101010101010101010101010101000111100110000111100001100111100,
64'b0011001111001100001100111100110011110000000011110000111111110000,
64'b1001100110011001011001100110011001011010101001011010010101011010,
64'b0011110011000011110000110011110010100101101001010101101001011010,
64'b0000000000000000000000000000000011111111000000001111111100000000,
64'b0011110011000011110000110011110010011001100110010110011001100110,
64'b0011110011000011110000110011110010101010101010101010101010101010,
64'b0000111111110000000011111111000000111100110000111100001100111100,
64'b1001011001101001011010011001011001011010010110100101101001011010,
64'b1100001100111100110000110011110000110011110011000011001111001100,
64'b1001100110011001011001100110011001011010101001011010010101011010,
64'b1010101010101010101010101010101000111100001111000011110000111100,
64'b0011110011000011110000110011110000111100110000111100001100111100,
64'b0110011001100110011001100110011011111111111111110000000000000000,
64'b0000111100001111111100001111000011111111111111110000000000000000,
64'b0011110000111100001111000011110001101001100101100110100110010110,
64'b0101101010100101101001010101101001101001011010011001011010010110,
64'b1010101010101010101010101010101010100101010110101010010101011010,
64'b0110011001100110011001100110011010101010010101010101010110101010,
64'b0011001100110011110011001100110000001111111100000000111111110000,
64'b0011001111001100001100111100110001101001100101100110100110010110,
64'b1100001100111100110000110011110001100110100110011001100101100110,
64'b1001100101100110100110010110011011001100110011001100110011001100,
64'b0011110000111100001111000011110011001100001100110011001111001100,
64'b0110011001100110011001100110011010100101010110101010010101011010,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b1001100101100110100110010110011010100101010110101010010101011010,
64'b1010101010101010101010101010101011111111000000001111111100000000,
64'b1010101001010101010101011010101010011001011001101001100101100110,
64'b0011110000111100001111000011110000110011001100111100110011001100,
64'b0110100110010110011010011001011010010110100101101001011010010110,
64'b0000000011111111111111110000000000110011001100111100110011001100,
64'b1001100101100110100110010110011010101010010101010101010110101010,
64'b0011110000111100001111000011110000111100110000111100001100111100,
64'b0000111111110000000011111111000011000011110000110011110000111100,
64'b0000000000000000000000000000000001011010010110100101101001011010,
64'b0000111111110000000011111111000000001111000011111111000011110000,
64'b0011110000111100001111000011110001100110100110011001100101100110,
64'b1001011001101001011010011001011011001100110011001100110011001100,
64'b1100110000110011001100111100110011001100001100110011001111001100,
64'b1001100101100110100110010110011011111111111111110000000000000000,
64'b0011110000111100001111000011110011000011110000110011110000111100,
64'b0101010101010101101010101010101011110000111100001111000011110000,
64'b1100110011001100110011001100110001101001100101100110100110010110,
64'b0101010101010101101010101010101011110000111100001111000011110000,
64'b0110100101101001100101101001011010011001100110010110011001100110,
64'b0000111111110000000011111111000001011010101001011010010101011010,
64'b0000000011111111111111110000000010100101010110101010010101011010,
64'b0000000000000000000000000000000010011001011001101001100101100110,
64'b0000000011111111111111110000000011111111000000001111111100000000,
64'b0000111111110000000011111111000001101001011010011001011010010110,
64'b0011110011000011110000110011110001011010010110100101101001011010,
64'b1010010110100101010110100101101000001111000011111111000011110000,
64'b0110100101101001100101101001011010101010101010101010101010101010,
64'b0000111111110000000011111111000010100101010110101010010101011010,
64'b1100110011001100110011001100110001010101101010100101010110101010,
64'b0101101001011010010110100101101011000011001111001100001100111100,
64'b1111000000001111000011111111000001101001011010011001011010010110,
64'b0000000000000000000000000000000001010101101010100101010110101010,
64'b0011001111001100001100111100110011111111000000001111111100000000,
64'b0000000000000000000000000000000010011001011001101001100101100110,
64'b0110100101101001100101101001011000000000000000000000000000000000,
64'b1111111111111111000000000000000011111111111111110000000000000000,
64'b1010101001010101010101011010101011000011001111001100001100111100,
64'b1010101010101010101010101010101011000011110000110011110000111100,
64'b1001011010010110100101101001011011110000111100001111000011110000,
64'b0011110000111100001111000011110000110011110011000011001111001100,
64'b1010010101011010101001010101101011000011001111001100001100111100,
64'b0000000011111111111111110000000011000011001111001100001100111100,
64'b0011110000111100001111000011110000000000000000000000000000000000,
64'b0011110000111100001111000011110001101001100101100110100110010110,
64'b1100001100111100110000110011110010011001100110010110011001100110,
64'b1001011010010110100101101001011011111111111111110000000000000000,
64'b1111111111111111000000000000000011000011110000110011110000111100,
64'b0000000011111111111111110000000000000000000000000000000000000000,
64'b1010101010101010101010101010101000000000000000000000000000000000,
64'b1001100110011001011001100110011001011010101001011010010101011010,
64'b0011110011000011110000110011110000001111111100000000111111110000,
64'b1100110011001100110011001100110001010101101010100101010110101010,
64'b0101101001011010010110100101101000001111000011111111000011110000,
64'b1100001100111100110000110011110011110000000011110000111111110000,
64'b0000111111110000000011111111000011110000000011110000111111110000,
64'b1010101010101010101010101010101000000000000000000000000000000000,
64'b0011001100110011110011001100110010010110011010010110100110010110,
64'b1001100110011001011001100110011000111100001111000011110000111100,
64'b0101101010100101101001010101101010101010101010101010101010101010,
64'b1111111111111111000000000000000010100101010110101010010101011010,
64'b1001011010010110100101101001011010101010101010101010101010101010,
64'b0110011001100110011001100110011000000000000000000000000000000000,
64'b0011110000111100001111000011110011001100001100110011001111001100,
64'b0000000000000000000000000000000010101010010101010101010110101010,
64'b0101010110101010010101011010101000110011001100111100110011001100,
64'b0110011001100110011001100110011011111111000000001111111100000000,
64'b1111111100000000111111110000000010101010010101010101010110101010,
64'b1111000011110000111100001111000010101010010101010101010110101010,
64'b1100001100111100110000110011110010101010101010101010101010101010,
64'b0101101001011010010110100101101010010110011010010110100110010110,
64'b1001011010010110100101101001011010100101010110101010010101011010,
64'b0110011010011001100110010110011011001100110011001100110011001100,
64'b1010101010101010101010101010101011001100001100110011001111001100,
64'b0110100110010110011010011001011011001100110011001100110011001100,
64'b0011110000111100001111000011110000000000000000000000000000000000,
64'b0000111111110000000011111111000000001111000011111111000011110000,
64'b0000000000000000000000000000000010011001100110010110011001100110,
64'b0011001100110011110011001100110001011010010110100101101001011010,
64'b0011110000111100001111000011110001010101010101011010101010101010,
64'b1111111111111111000000000000000000110011001100111100110011001100,
64'b1111111100000000111111110000000010011001100110010110011001100110,
64'b0000111111110000000011111111000001100110011001100110011001100110,
64'b0011001111001100001100111100110010010110011010010110100110010110,
64'b1100001100111100110000110011110001100110100110011001100101100110,
64'b1100001111000011001111000011110011110000111100001111000011110000,
64'b0110011001100110011001100110011000001111000011111111000011110000,
64'b0011110011000011110000110011110001011010010110100101101001011010,
64'b0000111111110000000011111111000000000000000000000000000000000000,
64'b0000000011111111111111110000000011111111000000001111111100000000,
64'b0000000000000000000000000000000010010110100101101001011010010110,
64'b1111000011110000111100001111000010011001011001101001100101100110,
64'b1010010101011010101001010101101011001100110011001100110011001100,
64'b0000000000000000000000000000000001011010010110100101101001011010,
64'b0101010101010101101010101010101010010110100101101001011010010110,
64'b1111111100000000111111110000000010010110100101101001011010010110,
64'b0000111100001111111100001111000010010110011010010110100110010110,
64'b1111000000001111000011111111000001101001011010011001011010010110,
64'b0000111111110000000011111111000001010101101010100101010110101010,
64'b1001011010010110100101101001011011111111000000001111111100000000,
64'b1111000000001111000011111111000010011001011001101001100101100110,
64'b1010101001010101010101011010101000000000000000000000000000000000,
64'b1111111111111111000000000000000011111111111111110000000000000000,
64'b1010101010101010101010101010101011000011001111001100001100111100,
64'b1111111100000000111111110000000011000011110000110011110000111100,
64'b1100110000110011001100111100110011110000111100001111000011110000,
64'b0000000000000000000000000000000000110011110011000011001111001100,
64'b1100110011001100110011001100110011000011001111001100001100111100,
64'b1010101010101010101010101010101011000011001111001100001100111100,
64'b1010101010101010101010101010101010010110011010010110100110010110,
64'b1111000011110000111100001111000001101001011010011001011010010110,
64'b0011001100110011110011001100110011000011001111001100001100111100,
64'b0101101010100101101001010101101001100110100110011001100101100110,
64'b1001011001101001011010011001011011111111111111110000000000000000,
64'b1010101010101010101010101010101001011010101001011010010101011010,
64'b1010010110100101010110100101101001101001100101100110100110010110,
64'b1100110000110011001100111100110000001111111100000000111111110000,
64'b0101010101010101101010101010101011111111111111110000000000000000,
64'b0110011010011001100110010110011011111111000000001111111100000000,
64'b0011110000111100001111000011110010100101101001010101101001011010,
64'b0110011010011001100110010110011010011001011001101001100101100110,
64'b1100110011001100110011001100110001101001100101100110100110010110,
64'b1100110011001100110011001100110010010110011010010110100110010110,
64'b0000111111110000000011111111000001101001100101100110100110010110,
64'b1100001111000011001111000011110001011010101001011010010101011010,
64'b0011110000111100001111000011110011000011110000110011110000111100,
64'b0000000000000000000000000000000010101010101010101010101010101010,
64'b1100110011001100110011001100110001100110100110011001100101100110,
64'b1001011001101001011010011001011010010110011010010110100110010110,
64'b0110100110010110011010011001011000000000111111111111111100000000,
64'b0011001100110011110011001100110000000000000000000000000000000000,
64'b0000111111110000000011111111000001010101010101011010101010101010,
64'b1001100101100110100110010110011000110011110011000011001111001100,
64'b1010010101011010101001010101101001101001011010011001011010010110,
64'b1001011010010110100101101001011011000011001111001100001100111100,
64'b0101101001011010010110100101101010010110011010010110100110010110,
64'b1111000000001111000011111111000010010110011010010110100110010110,
64'b0011110011000011110000110011110011001100001100110011001111001100,
64'b1111111111111111000000000000000010100101010110101010010101011010,
64'b1001011001101001011010011001011001100110011001100110011001100110,
64'b0101101001011010010110100101101011000011110000110011110000111100,
64'b1001100101100110100110010110011010010110011010010110100110010110,
64'b0101101001011010010110100101101001010101010101011010101010101010,
64'b1010010110100101010110100101101010101010101010101010101010101010,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b1111111111111111000000000000000010100101101001010101101001011010,
64'b1010101010101010101010101010101011000011001111001100001100111100,
64'b0000111111110000000011111111000010100101010110101010010101011010,
64'b0011001111001100001100111100110010010110011010010110100110010110,
64'b0000000011111111111111110000000010010110011010010110100110010110,
64'b0101101010100101101001010101101010100101101001010101101001011010,
64'b1010101010101010101010101010101001100110100110011001100101100110,
64'b1001011001101001011010011001011000111100001111000011110000111100,
64'b1001100101100110100110010110011000001111111100000000111111110000,
64'b1100001111000011001111000011110010010110011010010110100110010110,
64'b0011001111001100001100111100110001100110011001100110011001100110,
64'b0011001111001100001100111100110001100110011001100110011001100110,
64'b0101101001011010010110100101101011110000111100001111000011110000,
64'b0000000000000000000000000000000000110011110011000011001111001100,
64'b0110011001100110011001100110011001011010101001011010010101011010,
64'b1111111100000000111111110000000000110011110011000011001111001100,
64'b0000111100001111111100001111000000111100110000111100001100111100,
64'b0000111100001111111100001111000010010110011010010110100110010110,
64'b0101010110101010010101011010101010011001011001101001100101100110,
64'b0011110011000011110000110011110001101001011010011001011010010110,
64'b1010101010101010101010101010101010100101010110101010010101011010,
64'b1100001111000011001111000011110000000000111111111111111100000000,
64'b1010101001010101010101011010101000111100110000111100001100111100,
64'b0110100110010110011010011001011010010110100101101001011010010110,
64'b0101101001011010010110100101101000111100001111000011110000111100,
64'b0101010101010101101010101010101011111111000000001111111100000000,
64'b0011110000111100001111000011110000001111000011111111000011110000,
64'b0101101010100101101001010101101011001100001100110011001111001100,
64'b1100110011001100110011001100110001011010010110100101101001011010,
64'b0101010110101010010101011010101001011010101001011010010101011010,
64'b1010010101011010101001010101101010010110011010010110100110010110,
64'b1010101010101010101010101010101001101001011010011001011010010110,
64'b1010101010101010101010101010101011000011001111001100001100111100,
64'b1111000000001111000011111111000001100110100110011001100101100110,
64'b1010010101011010101001010101101011111111111111110000000000000000,
64'b0011110000111100001111000011110001011010101001011010010101011010,
64'b0101101001011010010110100101101001101001100101100110100110010110,
64'b0110011010011001100110010110011000001111111100000000111111110000,
64'b1010101001010101010101011010101011111111111111110000000000000000,
64'b1001100101100110100110010110011011111111000000001111111100000000,
64'b1010101010101010101010101010101010100101101001010101101001011010,
64'b1001011010010110100101101001011010011001011001101001100101100110,
64'b0011001100110011110011001100110011001100001100110011001111001100,
64'b1100110000110011001100111100110001100110100110011001100101100110,
64'b1100110011001100110011001100110001011010101001011010010101011010,
64'b1100110011001100110011001100110000000000000000000000000000000000,
64'b0000000011111111111111110000000001010101101010100101010110101010,
64'b0110011010011001100110010110011000000000000000000000000000000000,
64'b0000111111110000000011111111000011000011001111001100001100111100,
64'b0011001111001100001100111100110001011010010110100101101001011010,
64'b1100001111000011001111000011110001010101101010100101010110101010,
64'b1001100110011001011001100110011001100110100110011001100101100110,
64'b0110100101101001100101101001011001101001011010011001011010010110,
64'b1100110011001100110011001100110001010101010101011010101010101010,
64'b1100001100111100110000110011110001011010010110100101101001011010,
64'b0101101001011010010110100101101000001111000011111111000011110000,
64'b0101010101010101101010101010101010011001100110010110011001100110,
64'b0110100101101001100101101001011001010101101010100101010110101010,
64'b1010101001010101010101011010101011110000000011110000111111110000,
64'b0110100110010110011010011001011010100101010110101010010101011010,
64'b1100001111000011001111000011110010101010101010101010101010101010,
64'b0000111111110000000011111111000001010101101010100101010110101010,
64'b1100001100111100110000110011110011111111111111110000000000000000,
64'b0101101010100101101001010101101001100110011001100110011001100110,
64'b1111000000001111000011111111000010100101010110101010010101011010,
64'b0101010110101010010101011010101001010101101010100101010110101010,
64'b0011110011000011110000110011110000000000111111111111111100000000,
64'b1100001100111100110000110011110001010101101010100101010110101010,
64'b0011001111001100001100111100110011111111000000001111111100000000,
64'b0011110000111100001111000011110010010110100101101001011010010110,
64'b0101101010100101101001010101101010011001100110010110011001100110,
64'b1100001100111100110000110011110000000000111111111111111100000000,
64'b0000000000000000000000000000000001100110100110011001100101100110,
64'b1010010101011010101001010101101011001100110011001100110011001100,
64'b0000111111110000000011111111000000110011001100111100110011001100,
64'b0011110000111100001111000011110000000000000000000000000000000000,
64'b1001100101100110100110010110011010010110100101101001011010010110,
64'b1100110011001100110011001100110011001100001100110011001111001100,
64'b1010010110100101010110100101101000110011001100111100110011001100,
64'b1001011010010110100101101001011011111111111111110000000000000000,
64'b0110100110010110011010011001011001100110011001100110011001100110,
64'b0000111100001111111100001111000001010101010101011010101010101010,
64'b0000111111110000000011111111000011000011001111001100001100111100,
64'b1100110000110011001100111100110000111100001111000011110000111100,
64'b0101101010100101101001010101101001010101010101011010101010101010,
64'b0000000000000000000000000000000001101001011010011001011010010110,
64'b1100110000110011001100111100110001011010010110100101101001011010,
64'b0000000011111111111111110000000011110000111100001111000011110000,
64'b0000111111110000000011111111000010101010101010101010101010101010,
64'b1100001111000011001111000011110011000011001111001100001100111100,
64'b1111000011110000111100001111000000001111000011111111000011110000,
64'b0011001111001100001100111100110001011010010110100101101001011010,
64'b0110100110010110011010011001011010101010101010101010101010101010,
64'b1100001100111100110000110011110010010110100101101001011010010110,
64'b0101010110101010010101011010101011001100110011001100110011001100,
64'b0101101010100101101001010101101010101010010101010101010110101010,
64'b0011110000111100001111000011110000111100110000111100001100111100,
64'b0011110000111100001111000011110010010110011010010110100110010110,
64'b0011110011000011110000110011110011111111111111110000000000000000,
64'b1010010110100101010110100101101000110011110011000011001111001100,
64'b1111000011110000111100001111000001011010101001011010010101011010,
64'b0110011001100110011001100110011000000000111111111111111100000000,
64'b0101101010100101101001010101101010100101010110101010010101011010,
64'b0011001100110011110011001100110010011001100110010110011001100110,
64'b0011001100110011110011001100110010100101010110101010010101011010,
64'b0101101001011010010110100101101010101010010101010101010110101010,
64'b1100001100111100110000110011110000001111111100000000111111110000,
64'b1001100110011001011001100110011011110000111100001111000011110000,
64'b0011110011000011110000110011110000110011001100111100110011001100,
64'b1001011001101001011010011001011001011010101001011010010101011010,
64'b0101010101010101101010101010101010010110011010010110100110010110,
64'b0110011001100110011001100110011010101010101010101010101010101010,
64'b0011001111001100001100111100110010100101101001010101101001011010,
64'b1111000000001111000011111111000011001100001100110011001111001100,
64'b1111000000001111000011111111000001010101010101011010101010101010,
64'b1001100101100110100110010110011001100110100110011001100101100110,
64'b0011110011000011110000110011110000111100001111000011110000111100,
64'b0110011001100110011001100110011001100110100110011001100101100110,
64'b1111111111111111000000000000000000110011001100111100110011001100,
64'b1100001100111100110000110011110001010101101010100101010110101010,
64'b1001011010010110100101101001011011111111000000001111111100000000,
64'b1010101001010101010101011010101011110000111100001111000011110000,
64'b1010010101011010101001010101101001100110100110011001100101100110,
64'b0011110011000011110000110011110010010110011010010110100110010110,
64'b0000000011111111111111110000000001100110011001100110011001100110,
64'b1010010110100101010110100101101000110011110011000011001111001100,
64'b1010010101011010101001010101101010100101101001010101101001011010,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b0011110000111100001111000011110001101001011010011001011010010110,
64'b1001011010010110100101101001011010100101010110101010010101011010,
64'b1010101010101010101010101010101011000011110000110011110000111100,
64'b0110011010011001100110010110011001011010010110100101101001011010,
64'b0110100110010110011010011001011001100110011001100110011001100110,
64'b0110100110010110011010011001011011111111111111110000000000000000,
64'b0011001100110011110011001100110011111111000000001111111100000000,
64'b0110011010011001100110010110011011000011110000110011110000111100,
64'b1111000000001111000011111111000010010110011010010110100110010110,
64'b0101010101010101101010101010101010010110100101101001011010010110,
64'b1001100101100110100110010110011000001111000011111111000011110000,
64'b0110011010011001100110010110011000110011110011000011001111001100,
64'b0011110000111100001111000011110010010110100101101001011010010110,
64'b0000111111110000000011111111000011000011001111001100001100111100,
64'b1100001100111100110000110011110001100110100110011001100101100110,
64'b1100110011001100110011001100110000001111111100000000111111110000,
64'b1100001111000011001111000011110010011001011001101001100101100110,
64'b0110100110010110011010011001011000111100001111000011110000111100,
64'b1001011001101001011010011001011000000000000000000000000000000000,
64'b1111000011110000111100001111000001010101010101011010101010101010,
64'b0110100101101001100101101001011000001111111100000000111111110000,
64'b1010101001010101010101011010101010010110011010010110100110010110,
64'b0110011001100110011001100110011001101001100101100110100110010110,
64'b0110100101101001100101101001011011111111000000001111111100000000,
64'b1100001111000011001111000011110010100101101001010101101001011010,
64'b1010010101011010101001010101101011000011001111001100001100111100,
64'b0000000011111111111111110000000011110000000011110000111111110000,
64'b1111000000001111000011111111000011000011110000110011110000111100,
64'b1111000011110000111100001111000010101010010101010101010110101010,
64'b0000111111110000000011111111000011000011110000110011110000111100,
64'b0110100110010110011010011001011000001111111100000000111111110000,
64'b1001011001101001011010011001011000000000000000000000000000000000,
64'b0101010110101010010101011010101011001100110011001100110011001100,
64'b1100001100111100110000110011110010101010010101010101010110101010,
64'b1001100110011001011001100110011000111100110000111100001100111100,
64'b1001011010010110100101101001011010010110011010010110100110010110,
64'b1100001100111100110000110011110011111111111111110000000000000000,
64'b1010010101011010101001010101101000110011110011000011001111001100,
64'b0110011010011001100110010110011001011010101001011010010101011010,
64'b1111111111111111000000000000000000000000111111111111111100000000,
64'b1010101001010101010101011010101010100101010110101010010101011010,
64'b0101010110101010010101011010101010011001100110010110011001100110,
64'b0000000011111111111111110000000010100101010110101010010101011010,
64'b1100001100111100110000110011110001010101101010100101010110101010,
64'b1001100110011001011001100110011011110000000011110000111111110000,
64'b1001011001101001011010011001011011110000111100001111000011110000,
64'b1111111100000000111111110000000000001111000011111111000011110000,
64'b0000000011111111111111110000000000000000000000000000000000000000,
64'b1010010110100101010110100101101011001100001100110011001111001100,
64'b1001011010010110100101101001011001011010101001011010010101011010,
64'b1010101010101010101010101010101010100101101001010101101001011010,
64'b1100110011001100110011001100110011000011001111001100001100111100,
64'b0011110011000011110000110011110000001111000011111111000011110000,
64'b0000111100001111111100001111000010010110100101101001011010010110,
64'b0101101001011010010110100101101001010101101010100101010110101010,
64'b1010010101011010101001010101101001010101010101011010101010101010,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b1010010110100101010110100101101010101010010101010101010110101010,
64'b0000000000000000000000000000000001010101101010100101010110101010,
64'b1010101001010101010101011010101011111111000000001111111100000000,
64'b1111111100000000111111110000000010101010101010101010101010101010,
64'b0011110011000011110000110011110000001111000011111111000011110000,
64'b1111111100000000111111110000000001100110100110011001100101100110,
64'b0110011001100110011001100110011010011001011001101001100101100110,
64'b0011110000111100001111000011110001011010101001011010010101011010,
64'b1100110011001100110011001100110011111111000000001111111100000000,
64'b0101101010100101101001010101101001101001100101100110100110010110,
64'b1100001100111100110000110011110000110011001100111100110011001100,
64'b0110100101101001100101101001011011001100110011001100110011001100,
64'b0011110000111100001111000011110001011010010110100101101001011010,
64'b1010101001010101010101011010101010011001100110010110011001100110,
64'b0011110011000011110000110011110010011001100110010110011001100110,
64'b1100110000110011001100111100110011111111111111110000000000000000,
64'b0101010110101010010101011010101011001100110011001100110011001100,
64'b0101010110101010010101011010101011111111000000001111111100000000,
64'b1100001111000011001111000011110001101001011010011001011010010110,
64'b1001011010010110100101101001011001101001011010011001011010010110,
64'b1100001100111100110000110011110011001100001100110011001111001100,
64'b1100110000110011001100111100110001010101010101011010101010101010,
64'b1100001100111100110000110011110000111100110000111100001100111100,
64'b0000000011111111111111110000000011110000111100001111000011110000,
64'b0110011001100110011001100110011001011010010110100101101001011010,
64'b0110100110010110011010011001011000110011110011000011001111001100,
64'b1001100110011001011001100110011010010110100101101001011010010110,
64'b0101101010100101101001010101101010010110100101101001011010010110,
64'b1010010110100101010110100101101010101010101010101010101010101010,
64'b1001100110011001011001100110011001011010010110100101101001011010,
64'b0011001100110011110011001100110011111111111111110000000000000000,
64'b0000111111110000000011111111000011000011001111001100001100111100,
64'b0110100110010110011010011001011001101001100101100110100110010110,
64'b1111000000001111000011111111000010100101101001010101101001011010,
64'b0000111100001111111100001111000001100110011001100110011001100110,
64'b0101101010100101101001010101101001011010101001011010010101011010,
64'b1111111111111111000000000000000001010101101010100101010110101010,
64'b1001011010010110100101101001011000110011110011000011001111001100,
64'b1100001100111100110000110011110011110000111100001111000011110000,
64'b0000111100001111111100001111000001101001100101100110100110010110,
64'b1111000011110000111100001111000011000011001111001100001100111100,
64'b0110011001100110011001100110011011001100110011001100110011001100,
64'b1001011001101001011010011001011000110011110011000011001111001100,
64'b1111111111111111000000000000000000000000000000000000000000000000,
64'b0011110011000011110000110011110001011010101001011010010101011010,
64'b1001011001101001011010011001011000111100110000111100001100111100,
64'b1100110000110011001100111100110000110011110011000011001111001100,
64'b0110100101101001100101101001011010010110100101101001011010010110,
64'b0110100110010110011010011001011011001100001100110011001111001100,
64'b1111000011110000111100001111000010011001100110010110011001100110,
64'b1100110011001100110011001100110000001111000011111111000011110000,
64'b1100001100111100110000110011110011111111000000001111111100000000,
64'b0110011010011001100110010110011000111100110000111100001100111100,
64'b1100001111000011001111000011110011110000000011110000111111110000,
64'b1100001100111100110000110011110011110000111100001111000011110000,
64'b0011110000111100001111000011110000001111000011111111000011110000,
64'b0000111100001111111100001111000000000000000000000000000000000000,
64'b1100110000110011001100111100110011001100001100110011001111001100,
64'b0011110011000011110000110011110001011010101001011010010101011010,
64'b0110100101101001100101101001011010100101101001010101101001011010,
64'b0101010101010101101010101010101011000011001111001100001100111100,
64'b1001100101100110100110010110011000001111000011111111000011110000,
64'b1010010101011010101001010101101010010110100101101001011010010110,
64'b0101010110101010010101011010101001010101101010100101010110101010,
64'b1100001100111100110000110011110010101010101010101010101010101010,
64'b1100001111000011001111000011110011000011001111001100001100111100,
64'b1010010101011010101001010101101000111100001111000011110000111100,
64'b0101101010100101101001010101101010101010101010101010101010101010,
64'b0000111111110000000011111111000011111111111111110000000000000000,
64'b1111111100000000111111110000000000001111000011111111000011110000,
64'b1010010110100101010110100101101010011001100110010110011001100110,
64'b0101101010100101101001010101101011001100001100110011001111001100,
64'b0110100110010110011010011001011001010101101010100101010110101010,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b0110100101101001100101101001011011110000000011110000111111110000,
64'b1100110000110011001100111100110000110011110011000011001111001100,
64'b0011001100110011110011001100110010010110011010010110100110010110,
64'b0000111111110000000011111111000000000000000000000000000000000000,
64'b0011110011000011110000110011110001101001100101100110100110010110,
64'b1111000011110000111100001111000010011001100110010110011001100110,
64'b0011001100110011110011001100110000110011110011000011001111001100,
64'b1010101010101010101010101010101000000000111111111111111100000000,
64'b0101101001011010010110100101101011110000000011110000111111110000,
64'b1010010101011010101001010101101000000000000000000000000000000000,
64'b1100110000110011001100111100110000001111000011111111000011110000,
64'b0101101010100101101001010101101001010101010101011010101010101010,
64'b0000000011111111111111110000000000000000111111111111111100000000,
64'b1100110000110011001100111100110000001111111100000000111111110000,
64'b1111111111111111000000000000000011111111111111110000000000000000,
64'b1111111100000000111111110000000010011001100110010110011001100110,
64'b1001100101100110100110010110011001100110011001100110011001100110,
64'b1100001100111100110000110011110010010110011010010110100110010110,
64'b1100001111000011001111000011110000111100001111000011110000111100,
64'b0000111111110000000011111111000010100101101001010101101001011010,
64'b0110011010011001100110010110011011111111111111110000000000000000,
64'b1001011001101001011010011001011010101010010101010101010110101010,
64'b0101101010100101101001010101101010101010101010101010101010101010,
64'b1010010110100101010110100101101011111111000000001111111100000000,
64'b1010101001010101010101011010101001100110011001100110011001100110,
64'b0110100110010110011010011001011001010101010101011010101010101010,
64'b1010101010101010101010101010101010101010010101010101010110101010,
64'b1111000011110000111100001111000000000000000000000000000000000000,
64'b1111000000001111000011111111000010010110100101101001011010010110,
64'b1111000011110000111100001111000010010110100101101001011010010110,
64'b0101101010100101101001010101101000111100110000111100001100111100,
64'b0000111111110000000011111111000010100101010110101010010101011010,
64'b1010101001010101010101011010101000110011110011000011001111001100,
64'b1100001111000011001111000011110010101010101010101010101010101010,
64'b1001011001101001011010011001011010011001100110010110011001100110,
64'b0110011010011001100110010110011001100110011001100110011001100110,
64'b1001100101100110100110010110011011111111111111110000000000000000,
64'b1001100110011001011001100110011000111100001111000011110000111100,
64'b1001011001101001011010011001011011001100110011001100110011001100,
64'b1100110011001100110011001100110010011001100110010110011001100110,
64'b1111111100000000111111110000000010101010101010101010101010101010,
64'b0000000011111111111111110000000011000011001111001100001100111100,
64'b0101010110101010010101011010101011000011001111001100001100111100,
64'b1111111100000000111111110000000001101001100101100110100110010110,
64'b0011110000111100001111000011110011110000111100001111000011110000,
64'b1100110000110011001100111100110011110000000011110000111111110000,
64'b1010010110100101010110100101101011001100001100110011001111001100,
64'b0011001111001100001100111100110010011001100110010110011001100110,
64'b1111111111111111000000000000000000000000000000000000000000000000,
64'b1100001111000011001111000011110010101010101010101010101010101010,
64'b1111000011110000111100001111000001101001100101100110100110010110,
64'b1010101010101010101010101010101011001100001100110011001111001100,
64'b0101010101010101101010101010101000110011001100111100110011001100,
64'b1010010110100101010110100101101000111100001111000011110000111100,
64'b0101101010100101101001010101101001010101010101011010101010101010,
64'b1010101010101010101010101010101011000011001111001100001100111100,
64'b1100110011001100110011001100110010010110011010010110100110010110,
64'b1001100110011001011001100110011011111111000000001111111100000000,
64'b1111000000001111000011111111000000000000111111111111111100000000,
64'b1001100110011001011001100110011010100101101001010101101001011010,
64'b0000000000000000000000000000000010010110100101101001011010010110,
64'b1001011010010110100101101001011010101010101010101010101010101010,
64'b0000111111110000000011111111000011001100110011001100110011001100,
64'b1001100101100110100110010110011000111100110000111100001100111100,
64'b1111000000001111000011111111000000001111000011111111000011110000,
64'b1100001111000011001111000011110001011010010110100101101001011010,
64'b1100001100111100110000110011110010100101010110101010010101011010,
64'b1100001111000011001111000011110011001100110011001100110011001100,
64'b1010101010101010101010101010101010100101010110101010010101011010,
64'b1100001111000011001111000011110010010110011010010110100110010110,
64'b1010101001010101010101011010101001010101010101011010101010101010,
64'b0101010101010101101010101010101011111111111111110000000000000000,
64'b1001011001101001011010011001011010011001011001101001100101100110,
64'b0000111100001111111100001111000001101001100101100110100110010110,
64'b0101010110101010010101011010101011001100110011001100110011001100,
64'b1010101001010101010101011010101011110000111100001111000011110000,
64'b0000111100001111111100001111000011110000000011110000111111110000,
64'b0011110000111100001111000011110001010101101010100101010110101010,
64'b1010101001010101010101011010101010011001011001101001100101100110,
64'b0000000011111111111111110000000011001100001100110011001111001100,
64'b1010101010101010101010101010101011110000111100001111000011110000,
64'b1010101010101010101010101010101000110011110011000011001111001100,
64'b1010010101011010101001010101101000111100110000111100001100111100,
64'b1001100110011001011001100110011001100110011001100110011001100110,
64'b0110011001100110011001100110011010101010101010101010101010101010,
64'b1001011001101001011010011001011001101001011010011001011010010110,
64'b0101010110101010010101011010101000111100110000111100001100111100,
64'b1001100110011001011001100110011011110000111100001111000011110000,
64'b0011001100110011110011001100110011111111000000001111111100000000,
64'b0101010110101010010101011010101000000000111111111111111100000000,
64'b1010010101011010101001010101101010011001100110010110011001100110,
64'b0011001100110011110011001100110011000011110000110011110000111100,
64'b0101010101010101101010101010101000001111000011111111000011110000,
64'b0110011001100110011001100110011001010101101010100101010110101010,
64'b1100110011001100110011001100110011110000111100001111000011110000,
64'b0110011010011001100110010110011011110000000011110000111111110000,
64'b0011110000111100001111000011110010010110100101101001011010010110,
64'b1001011010010110100101101001011011001100110011001100110011001100,
64'b0011110011000011110000110011110011000011001111001100001100111100,
64'b1001100110011001011001100110011001011010101001011010010101011010,
64'b0011110000111100001111000011110001010101101010100101010110101010,
64'b0101101001011010010110100101101011111111111111110000000000000000,
64'b1001100110011001011001100110011011111111111111110000000000000000,
64'b1100110000110011001100111100110010010110100101101001011010010110,
64'b1111000011110000111100001111000010100101010110101010010101011010,
64'b0110011001100110011001100110011001010101101010100101010110101010,
64'b1001011010010110100101101001011010011001100110010110011001100110,
64'b1111000011110000111100001111000011111111000000001111111100000000,
64'b0110100101101001100101101001011010101010010101010101010110101010,
64'b1010010101011010101001010101101001101001100101100110100110010110,
64'b1100001100111100110000110011110011110000111100001111000011110000,
64'b1111000000001111000011111111000011110000000011110000111111110000,
64'b1001011010010110100101101001011011001100001100110011001111001100,
64'b1010010101011010101001010101101010011001100110010110011001100110,
64'b0011001111001100001100111100110000000000000000000000000000000000,
64'b0011110000111100001111000011110010101010101010101010101010101010,
64'b1010010110100101010110100101101001101001100101100110100110010110,
64'b0101010110101010010101011010101011001100001100110011001111001100,
64'b0011110000111100001111000011110000110011001100111100110011001100,
64'b1100001100111100110000110011110000111100001111000011110000111100,
64'b1111111100000000111111110000000010101010101010101010101010101010,
64'b1100110000110011001100111100110001100110100110011001100101100110,
64'b0110100101101001100101101001011011000011001111001100001100111100,
64'b1100110011001100110011001100110010101010101010101010101010101010,
64'b0110100110010110011010011001011011110000111100001111000011110000,
64'b1111111111111111000000000000000010011001100110010110011001100110,
64'b0011001111001100001100111100110011001100110011001100110011001100,
64'b0101101001011010010110100101101011110000111100001111000011110000,
64'b1001100110011001011001100110011011000011110000110011110000111100,
64'b0000111100001111111100001111000011000011110000110011110000111100,
64'b0110011010011001100110010110011000111100001111000011110000111100,
64'b1010010110100101010110100101101011110000111100001111000011110000,
64'b0000000000000000000000000000000010101010010101010101010110101010,
64'b0110011001100110011001100110011000000000000000000000000000000000,
64'b1100001100111100110000110011110011000011110000110011110000111100,
64'b0000000011111111111111110000000001011010101001011010010101011010,
64'b1001011010010110100101101001011011001100110011001100110011001100,
64'b0101010101010101101010101010101011111111000000001111111100000000,
64'b1111111111111111000000000000000000111100001111000011110000111100,
64'b1001011001101001011010011001011001011010010110100101101001011010,
64'b0110100110010110011010011001011011111111000000001111111100000000,
64'b1010010110100101010110100101101000001111111100000000111111110000,
64'b0101101010100101101001010101101010100101010110101010010101011010,
64'b0000111111110000000011111111000010100101010110101010010101011010,
64'b0011110011000011110000110011110011111111000000001111111100000000,
64'b1010101010101010101010101010101000110011001100111100110011001100,
64'b0101101001011010010110100101101010101010101010101010101010101010,
64'b0011110000111100001111000011110000001111111100000000111111110000,
64'b1001011010010110100101101001011001100110100110011001100101100110,
64'b1010010101011010101001010101101001011010010110100101101001011010,
64'b1010010101011010101001010101101011111111111111110000000000000000,
64'b0101010101010101101010101010101000001111111100000000111111110000,
64'b1010010110100101010110100101101000110011110011000011001111001100,
64'b1100110000110011001100111100110011111111111111110000000000000000,
64'b1010101001010101010101011010101000000000111111111111111100000000,
64'b0110100110010110011010011001011011001100001100110011001111001100,
64'b1100110011001100110011001100110011001100001100110011001111001100,
64'b0101010110101010010101011010101011111111111111110000000000000000,
64'b0110011001100110011001100110011011110000111100001111000011110000,
64'b0101010110101010010101011010101001100110011001100110011001100110,
64'b1010010101011010101001010101101010101010010101010101010110101010,
64'b1100001100111100110000110011110011000011110000110011110000111100,
64'b1100110000110011001100111100110010011001011001101001100101100110,
64'b1100110000110011001100111100110000000000000000000000000000000000,
64'b1100110011001100110011001100110010101010010101010101010110101010,
64'b1001100101100110100110010110011000001111000011111111000011110000,
64'b1010010110100101010110100101101000000000000000000000000000000000,
64'b1001100110011001011001100110011001010101010101011010101010101010,
64'b1001011001101001011010011001011010100101101001010101101001011010,
64'b1111000011110000111100001111000010100101101001010101101001011010,
64'b0011001100110011110011001100110010101010101010101010101010101010,
64'b0011110000111100001111000011110001010101101010100101010110101010,
64'b1100110011001100110011001100110000111100001111000011110000111100,
64'b1010101010101010101010101010101000110011001100111100110011001100,
64'b1001100101100110100110010110011010100101010110101010010101011010,
64'b1100001111000011001111000011110001101001011010011001011010010110,
64'b1100110000110011001100111100110000000000000000000000000000000000,
64'b1010010110100101010110100101101000110011001100111100110011001100,
64'b1111000000001111000011111111000001010101101010100101010110101010,
64'b0110100110010110011010011001011010101010101010101010101010101010,
64'b0000111100001111111100001111000011001100110011001100110011001100,
64'b1001100101100110100110010110011010011001011001101001100101100110,
64'b0011001100110011110011001100110010011001011001101001100101100110,
64'b0101010101010101101010101010101001100110011001100110011001100110,
64'b1010010101011010101001010101101000110011001100111100110011001100,
64'b1001011010010110100101101001011000001111111100000000111111110000,
64'b1010101001010101010101011010101001011010010110100101101001011010,
64'b1010101010101010101010101010101001100110100110011001100101100110,
64'b1100001100111100110000110011110011000011001111001100001100111100,
64'b1100110000110011001100111100110010101010101010101010101010101010,
64'b0110011010011001100110010110011011110000111100001111000011110000,
64'b1001100110011001011001100110011010011001100110010110011001100110,
64'b1100110000110011001100111100110011001100110011001100110011001100,
64'b0110011010011001100110010110011011110000111100001111000011110000,
64'b0110011001100110011001100110011011000011110000110011110000111100,
64'b1001011001101001011010011001011011000011110000110011110000111100,
64'b1100001111000011001111000011110000111100001111000011110000111100,
64'b0110011010011001100110010110011011110000111100001111000011110000,
64'b1010010101011010101001010101101001010101101010100101010110101010,
64'b1001100110011001011001100110011011111111111111110000000000000000,
64'b0110011001100110011001100110011010101010101010101010101010101010,
64'b1111000000001111000011111111000010010110011010010110100110010110,
64'b0000111100001111111100001111000010100101010110101010010101011010,
64'b0110100101101001100101101001011000000000111111111111111100000000,
64'b1001011010010110100101101001011000001111111100000000111111110000,
64'b1010010110100101010110100101101000000000000000000000000000000000,
64'b0110100101101001100101101001011001100110100110011001100101100110,
64'b1001011010010110100101101001011000000000111111111111111100000000,
64'b0011110011000011110000110011110011000011110000110011110000111100,
64'b1010010101011010101001010101101000000000111111111111111100000000,
64'b0110100101101001100101101001011011111111000000001111111100000000,
64'b1001100101100110100110010110011010101010101010101010101010101010,
64'b0101101010100101101001010101101011001100001100110011001111001100,
64'b1111111111111111000000000000000000001111000011111111000011110000,
64'b1100110000110011001100111100110011110000000011110000111111110000,
64'b0011110000111100001111000011110000001111000011111111000011110000,
64'b1001011001101001011010011001011000000000000000000000000000000000,
64'b0101101001011010010110100101101010011001100110010110011001100110,
64'b0110100110010110011010011001011001011010010110100101101001011010,
64'b1111000000001111000011111111000001011010010110100101101001011010,
64'b0110011010011001100110010110011001011010010110100101101001011010,
64'b1001011010010110100101101001011011000011110000110011110000111100,
64'b1100001100111100110000110011110011110000111100001111000011110000,
64'b1100001100111100110000110011110001010101010101011010101010101010,
64'b1111000011110000111100001111000010101010101010101010101010101010,
64'b1010101010101010101010101010101000001111000011111111000011110000,
64'b1100001111000011001111000011110001010101101010100101010110101010,
64'b0110100101101001100101101001011010101010010101010101010110101010,
64'b1100110011001100110011001100110001010101101010100101010110101010,
64'b1100001100111100110000110011110010101010101010101010101010101010,
64'b1010101010101010101010101010101000111100001111000011110000111100,
64'b0110011010011001100110010110011010011001011001101001100101100110,
64'b1001100101100110100110010110011000110011110011000011001111001100,
64'b0110011001100110011001100110011000110011110011000011001111001100,
64'b0000111100001111111100001111000000001111111100000000111111110000,
64'b0101010110101010010101011010101001010101101010100101010110101010,
64'b1111000000001111000011111111000011001100110011001100110011001100,
64'b1001100101100110100110010110011001100110011001100110011001100110,
64'b1100110011001100110011001100110011111111000000001111111100000000,
64'b0000111111110000000011111111000010011001100110010110011001100110,
64'b0110100110010110011010011001011000110011001100111100110011001100,
64'b0101101001011010010110100101101010011001100110010110011001100110,
64'b1111000000001111000011111111000011001100110011001100110011001100,
64'b1100110011001100110011001100110000001111111100000000111111110000,
64'b1100001111000011001111000011110011000011110000110011110000111100,
64'b0110100101101001100101101001011000001111000011111111000011110000,
64'b0011110000111100001111000011110000001111000011111111000011110000,
64'b1111111100000000111111110000000000000000111111111111111100000000,
64'b1001100110011001011001100110011000110011001100111100110011001100,
64'b0000000011111111111111110000000011110000111100001111000011110000,
64'b1001011010010110100101101001011000111100001111000011110000111100,
64'b1001011001101001011010011001011010011001011001101001100101100110,
64'b0110100110010110011010011001011001010101010101011010101010101010,
64'b1111000000001111000011111111000010010110100101101001011010010110,
64'b0101101001011010010110100101101011111111000000001111111100000000,
64'b1111111100000000111111110000000010100101101001010101101001011010,
64'b0110100110010110011010011001011000110011001100111100110011001100,
64'b0101010110101010010101011010101001010101101010100101010110101010,
64'b1111000000001111000011111111000011001100001100110011001111001100,
64'b1010101001010101010101011010101001011010101001011010010101011010,
64'b1001100101100110100110010110011000110011110011000011001111001100,
64'b1001100110011001011001100110011011111111111111110000000000000000,
64'b0101010101010101101010101010101001010101101010100101010110101010,
64'b0000111111110000000011111111000001101001100101100110100110010110,
64'b1111000011110000111100001111000001101001011010011001011010010110,
64'b1111111100000000111111110000000011001100110011001100110011001100,
64'b1100110000110011001100111100110001101001100101100110100110010110,
64'b1111000011110000111100001111000011111111111111110000000000000000,
64'b0000000000000000000000000000000000110011110011000011001111001100,
64'b0000111100001111111100001111000001011010010110100101101001011010,
64'b0110100101101001100101101001011010011001100110010110011001100110,
64'b1001100101100110100110010110011000001111000011111111000011110000,
64'b1001011010010110100101101001011001100110100110011001100101100110,
64'b0000111111110000000011111111000010100101101001010101101001011010,
64'b1001100110011001011001100110011000000000000000000000000000000000,
64'b0110011001100110011001100110011010011001100110010110011001100110,
64'b0011001111001100001100111100110011000011001111001100001100111100,
64'b0011001100110011110011001100110001101001100101100110100110010110,
64'b1001011010010110100101101001011001011010010110100101101001011010,
64'b1100001111000011001111000011110000111100110000111100001100111100,
64'b0011110000111100001111000011110000000000000000000000000000000000,
64'b1111111111111111000000000000000010100101101001010101101001011010,
64'b1100110011001100110011001100110000110011110011000011001111001100,
64'b0011001111001100001100111100110000111100001111000011110000111100,
64'b1111000011110000111100001111000001010101101010100101010110101010,
64'b1100110000110011001100111100110001101001011010011001011010010110,
64'b0110011001100110011001100110011010011001011001101001100101100110,
64'b1001100110011001011001100110011010101010101010101010101010101010,
64'b1001011010010110100101101001011000111100001111000011110000111100,
64'b1001011010010110100101101001011010100101010110101010010101011010,
64'b1111000011110000111100001111000010010110011010010110100110010110,
64'b0110100110010110011010011001011000110011110011000011001111001100,
64'b0000111111110000000011111111000011110000000011110000111111110000,
64'b1010010101011010101001010101101010101010101010101010101010101010,
64'b0000000000000000000000000000000000110011110011000011001111001100,
64'b0101101001011010010110100101101010100101101001010101101001011010,
64'b0000111100001111111100001111000000001111111100000000111111110000,
64'b1111111100000000111111110000000000110011001100111100110011001100,
64'b0000111100001111111100001111000011000011001111001100001100111100,
64'b1001011010010110100101101001011001101001011010011001011010010110,
64'b0011110000111100001111000011110011001100110011001100110011001100,
64'b0110100110010110011010011001011000001111111100000000111111110000,
64'b1100001100111100110000110011110000110011110011000011001111001100,
64'b1111111100000000111111110000000000111100110000111100001100111100,
64'b0011110011000011110000110011110010100101101001010101101001011010,
64'b0000000011111111111111110000000000000000111111111111111100000000,
64'b1100110000110011001100111100110001100110011001100110011001100110,
64'b0000000000000000000000000000000000001111000011111111000011110000,
64'b0011001111001100001100111100110000110011110011000011001111001100,
64'b1111111100000000111111110000000010101010010101010101010110101010,
64'b0101010101010101101010101010101011110000111100001111000011110000,
64'b1111111100000000111111110000000001011010101001011010010101011010,
64'b0110100110010110011010011001011011000011001111001100001100111100,
64'b0000111111110000000011111111000001011010010110100101101001011010,
64'b0011110011000011110000110011110000000000111111111111111100000000,
64'b0000111111110000000011111111000011110000111100001111000011110000,
64'b1111111111111111000000000000000001011010101001011010010101011010,
64'b1111000000001111000011111111000010011001011001101001100101100110,
64'b0101010101010101101010101010101001010101010101011010101010101010,
64'b1010010110100101010110100101101010010110100101101001011010010110,
64'b1010101010101010101010101010101011111111000000001111111100000000,
64'b0000111100001111111100001111000010100101101001010101101001011010,
64'b1111111111111111000000000000000000110011001100111100110011001100,
64'b1100110011001100110011001100110001010101101010100101010110101010,
64'b0101010101010101101010101010101011001100001100110011001111001100,
64'b0011110011000011110000110011110001011010101001011010010101011010,
64'b0000000011111111111111110000000000110011110011000011001111001100,
64'b1111000000001111000011111111000011111111111111110000000000000000,
64'b0101010110101010010101011010101001010101101010100101010110101010,
64'b0101101010100101101001010101101011001100001100110011001111001100,
64'b1001100101100110100110010110011010010110011010010110100110010110,
64'b0110100101101001100101101001011011111111000000001111111100000000,
64'b1111000011110000111100001111000000000000111111111111111100000000,
64'b0011001111001100001100111100110001010101010101011010101010101010,
64'b0110011001100110011001100110011000110011001100111100110011001100,
64'b0101010110101010010101011010101010101010101010101010101010101010,
64'b0110011001100110011001100110011010100101101001010101101001011010,
64'b0011110011000011110000110011110011000011110000110011110000111100,
64'b0101101010100101101001010101101010100101101001010101101001011010,
64'b1111111111111111000000000000000011111111000000001111111100000000,
64'b1001011001101001011010011001011011000011001111001100001100111100,
64'b0000111111110000000011111111000010100101010110101010010101011010,
64'b1001011010010110100101101001011000001111000011111111000011110000,
64'b1111000000001111000011111111000010010110011010010110100110010110,
64'b1010101001010101010101011010101001010101010101011010101010101010,
64'b1010010101011010101001010101101011111111111111110000000000000000,
64'b0011110011000011110000110011110001100110011001100110011001100110,
64'b0101101001011010010110100101101001011010010110100101101001011010,
64'b0110011010011001100110010110011001100110011001100110011001100110,
64'b0101101001011010010110100101101000110011110011000011001111001100,
64'b1100110011001100110011001100110010100101010110101010010101011010,
64'b0011110000111100001111000011110010011001011001101001100101100110,
64'b0101010101010101101010101010101001010101010101011010101010101010,
64'b0000000000000000000000000000000011110000000011110000111111110000,
64'b0101101001011010010110100101101000110011110011000011001111001100,
64'b1001100110011001011001100110011011111111000000001111111100000000,
64'b1001100110011001011001100110011010010110011010010110100110010110,
64'b1111000011110000111100001111000001100110011001100110011001100110,
64'b1001011001101001011010011001011010101010101010101010101010101010,
64'b1100001111000011001111000011110010010110100101101001011010010110,
64'b1111111100000000111111110000000000110011110011000011001111001100,
64'b1001011001101001011010011001011000111100001111000011110000111100,
64'b1111111100000000111111110000000000001111000011111111000011110000,
64'b1100110000110011001100111100110011001100001100110011001111001100,
64'b0101010101010101101010101010101011000011110000110011110000111100,
64'b0011001100110011110011001100110011001100110011001100110011001100,
64'b0011110011000011110000110011110010101010010101010101010110101010,
64'b0011110000111100001111000011110001011010010110100101101001011010,
64'b1001011010010110100101101001011011111111111111110000000000000000,
64'b1001011010010110100101101001011000111100110000111100001100111100,
64'b0101010110101010010101011010101010010110100101101001011010010110,
64'b0011110011000011110000110011110011001100110011001100110011001100,
64'b1010010101011010101001010101101011000011001111001100001100111100,
64'b0101010101010101101010101010101000001111000011111111000011110000,
64'b0011110011000011110000110011110000001111111100000000111111110000,
64'b0101010101010101101010101010101011111111000000001111111100000000,
64'b0000111100001111111100001111000010100101101001010101101001011010,
64'b0110011001100110011001100110011010100101010110101010010101011010,
64'b0101101001011010010110100101101001011010010110100101101001011010,
64'b0101101010100101101001010101101000110011001100111100110011001100,
64'b1010010101011010101001010101101010011001011001101001100101100110,
64'b1001100110011001011001100110011000000000000000000000000000000000,
64'b0101101001011010010110100101101001011010101001011010010101011010,
64'b0101101001011010010110100101101001101001100101100110100110010110,
64'b0000000011111111111111110000000011110000111100001111000011110000,
64'b0101010101010101101010101010101011110000000011110000111111110000,
64'b1010101010101010101010101010101011111111000000001111111100000000,
64'b0000111100001111111100001111000010101010010101010101010110101010,
64'b0000000000000000000000000000000011111111111111110000000000000000,
64'b0110100101101001100101101001011000110011110011000011001111001100,
64'b1100110000110011001100111100110001100110100110011001100101100110,
64'b1100110000110011001100111100110000110011110011000011001111001100,
64'b0101101001011010010110100101101011110000111100001111000011110000,
64'b1001011010010110100101101001011010010110100101101001011010010110,
64'b0110011010011001100110010110011010101010101010101010101010101010,
64'b0000000000000000000000000000000011001100001100110011001111001100,
64'b0101101010100101101001010101101010010110011010010110100110010110,
64'b0000111100001111111100001111000011111111000000001111111100000000,
64'b0101010110101010010101011010101000000000111111111111111100000000,
64'b0000000000000000000000000000000001010101010101011010101010101010,
64'b1010101010101010101010101010101000110011001100111100110011001100,
64'b1100110011001100110011001100110010101010101010101010101010101010,
64'b1111111111111111000000000000000010100101101001010101101001011010,
64'b1111111100000000111111110000000011000011110000110011110000111100,
64'b0101101001011010010110100101101010100101101001010101101001011010,
64'b0000111100001111111100001111000011111111000000001111111100000000,
64'b1100110011001100110011001100110011000011001111001100001100111100,
64'b0110100101101001100101101001011000111100110000111100001100111100,
64'b1010101010101010101010101010101010010110011010010110100110010110,
64'b1100110000110011001100111100110011111111000000001111111100000000,
64'b0101010110101010010101011010101010100101101001010101101001011010,
64'b1001100110011001011001100110011011001100001100110011001111001100,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1100110011001100110011001100110000001111111100000000111111110000,
64'b1111000011110000111100001111000000000000000000000000000000000000,
64'b0000000000000000000000000000000000001111000011111111000011110000,
64'b0101010101010101101010101010101011111111111111110000000000000000,
64'b0011001111001100001100111100110001100110100110011001100101100110,
64'b1111111100000000111111110000000011000011001111001100001100111100,
64'b0101101001011010010110100101101000000000000000000000000000000000,
64'b0011001100110011110011001100110010101010101010101010101010101010,
64'b1111111100000000111111110000000000001111000011111111000011110000,
64'b0110011001100110011001100110011000111100001111000011110000111100,
64'b0110100101101001100101101001011011000011001111001100001100111100,
64'b0000111111110000000011111111000010010110011010010110100110010110,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b1010010101011010101001010101101001010101010101011010101010101010,
64'b1001100101100110100110010110011001100110011001100110011001100110,
64'b0011110011000011110000110011110011000011110000110011110000111100,
64'b1001011001101001011010011001011011110000000011110000111111110000,
64'b0101101001011010010110100101101010010110100101101001011010010110,
64'b0110100110010110011010011001011011001100110011001100110011001100,
64'b0011110000111100001111000011110000001111111100000000111111110000,
64'b1010101001010101010101011010101011001100110011001100110011001100,
64'b1100110000110011001100111100110011111111000000001111111100000000,
64'b0101010101010101101010101010101010100101010110101010010101011010,
64'b0011001111001100001100111100110011110000000011110000111111110000,
64'b1001100110011001011001100110011000111100110000111100001100111100,
64'b1001011010010110100101101001011001011010010110100101101001011010,
64'b1001100110011001011001100110011011001100110011001100110011001100,
64'b1010010110100101010110100101101010010110100101101001011010010110,
64'b1100110011001100110011001100110000001111111100000000111111110000,
64'b1100110011001100110011001100110010101010010101010101010110101010,
64'b0110011010011001100110010110011001101001100101100110100110010110,
64'b1010101010101010101010101010101011110000111100001111000011110000,
64'b0000000000000000000000000000000011111111000000001111111100000000,
64'b1001100110011001011001100110011011110000111100001111000011110000,
64'b1010010110100101010110100101101011111111111111110000000000000000,
64'b0110011001100110011001100110011011001100001100110011001111001100,
64'b1010010110100101010110100101101000000000111111111111111100000000,
64'b0011110000111100001111000011110001011010101001011010010101011010,
64'b0110100110010110011010011001011010011001011001101001100101100110,
64'b0011110000111100001111000011110011110000111100001111000011110000,
64'b1001100101100110100110010110011011000011001111001100001100111100,
64'b0101101001011010010110100101101000000000111111111111111100000000,
64'b1111000011110000111100001111000000110011001100111100110011001100,
64'b1100001111000011001111000011110010010110011010010110100110010110,
64'b0110011001100110011001100110011011111111000000001111111100000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0110011010011001100110010110011010100101101001010101101001011010,
64'b0000000000000000000000000000000010011001011001101001100101100110,
64'b1111111111111111000000000000000011001100110011001100110011001100,
64'b1100001100111100110000110011110010100101101001010101101001011010,
64'b1001011010010110100101101001011001010101010101011010101010101010,
64'b0101101010100101101001010101101000001111000011111111000011110000,
64'b0101101001011010010110100101101010101010101010101010101010101010,
64'b1010010110100101010110100101101010010110011010010110100110010110,
64'b0000111100001111111100001111000011000011001111001100001100111100,
64'b1010010110100101010110100101101000000000111111111111111100000000,
64'b1111000000001111000011111111000001101001100101100110100110010110,
64'b0000000011111111111111110000000011000011001111001100001100111100,
64'b0000111111110000000011111111000000001111111100000000111111110000,
64'b0011001111001100001100111100110010011001011001101001100101100110,
64'b0011001111001100001100111100110001101001011010011001011010010110,
64'b0110100101101001100101101001011011110000111100001111000011110000,
64'b1010101001010101010101011010101000110011110011000011001111001100,
64'b1111000011110000111100001111000001100110011001100110011001100110,
64'b1010101001010101010101011010101001010101101010100101010110101010,
64'b1100110011001100110011001100110001100110011001100110011001100110,
64'b0101010110101010010101011010101000111100110000111100001100111100,
64'b0110100101101001100101101001011001011010101001011010010101011010,
64'b1100001111000011001111000011110011111111111111110000000000000000,
64'b0101010110101010010101011010101010010110011010010110100110010110,
64'b1100001100111100110000110011110011110000000011110000111111110000,
64'b0101101001011010010110100101101011111111000000001111111100000000,
64'b1111111100000000111111110000000001101001011010011001011010010110,
64'b1001011001101001011010011001011011000011001111001100001100111100,
64'b1010101001010101010101011010101001010101101010100101010110101010,
64'b0110100101101001100101101001011000001111000011111111000011110000,
64'b0110011001100110011001100110011000111100001111000011110000111100,
64'b0101010101010101101010101010101000110011001100111100110011001100,
64'b0000111111110000000011111111000000111100001111000011110000111100,
64'b0101010101010101101010101010101011110000000011110000111111110000,
64'b1111111111111111000000000000000001100110100110011001100101100110,
64'b1111111111111111000000000000000010101010101010101010101010101010,
64'b0110011001100110011001100110011010010110011010010110100110010110,
64'b0110011001100110011001100110011010101010010101010101010110101010,
64'b0011110000111100001111000011110010101010101010101010101010101010,
64'b1111111111111111000000000000000001101001100101100110100110010110,
64'b0011110011000011110000110011110001011010101001011010010101011010,
64'b1001100110011001011001100110011000110011001100111100110011001100,
64'b0110100110010110011010011001011011111111000000001111111100000000,
64'b1001011010010110100101101001011010100101010110101010010101011010,
64'b1100110011001100110011001100110011110000111100001111000011110000,
64'b1010101001010101010101011010101010100101010110101010010101011010,
64'b1100110011001100110011001100110000000000111111111111111100000000,
64'b1010101010101010101010101010101001101001011010011001011010010110,
64'b1010101010101010101010101010101001100110011001100110011001100110,
64'b1001011010010110100101101001011000111100110000111100001100111100,
64'b0011110000111100001111000011110010011001100110010110011001100110,
64'b0000111111110000000011111111000001100110011001100110011001100110,
64'b1010101010101010101010101010101010010110011010010110100110010110,
64'b0101101010100101101001010101101011001100001100110011001111001100,
64'b1001011010010110100101101001011001011010010110100101101001011010,
64'b1001011001101001011010011001011001010101010101011010101010101010,
64'b1100001100111100110000110011110011001100001100110011001111001100,
64'b1111000011110000111100001111000011111111000000001111111100000000,
64'b0011001100110011110011001100110011001100001100110011001111001100,
64'b0101101001011010010110100101101011111111111111110000000000000000,
64'b1100110011001100110011001100110001101001100101100110100110010110,
64'b1100110011001100110011001100110010010110100101101001011010010110,
64'b1100001100111100110000110011110011110000000011110000111111110000,
64'b0000111111110000000011111111000010010110100101101001011010010110,
64'b1111111100000000111111110000000010010110100101101001011010010110,
64'b0110011001100110011001100110011000111100110000111100001100111100,
64'b1100110000110011001100111100110010100101101001010101101001011010,
64'b0110100110010110011010011001011010011001011001101001100101100110,
64'b0011110011000011110000110011110011001100110011001100110011001100,
64'b0101101010100101101001010101101010100101101001010101101001011010,
64'b1111111100000000111111110000000001010101010101011010101010101010,
64'b1111000011110000111100001111000000001111000011111111000011110000,
64'b1001100101100110100110010110011010101010101010101010101010101010,
64'b1111000011110000111100001111000010010110011010010110100110010110,
64'b1111000011110000111100001111000011000011001111001100001100111100,
64'b1111000000001111000011111111000000000000111111111111111100000000,
64'b0000000011111111111111110000000001101001100101100110100110010110,
64'b0000000000000000000000000000000011000011001111001100001100111100,
64'b0101010101010101101010101010101010010110100101101001011010010110,
64'b1001011001101001011010011001011010100101010110101010010101011010,
64'b0110011001100110011001100110011000110011110011000011001111001100,
64'b1111111100000000111111110000000000111100001111000011110000111100,
64'b1111111100000000111111110000000011001100110011001100110011001100,
64'b1111111100000000111111110000000010010110100101101001011010010110,
64'b1111111111111111000000000000000010010110100101101001011010010110,
64'b1111111100000000111111110000000001100110100110011001100101100110,
64'b1001011010010110100101101001011001100110100110011001100101100110,
64'b1111000000001111000011111111000010011001100110010110011001100110,
64'b0011001111001100001100111100110011110000000011110000111111110000,
64'b1111111111111111000000000000000001010101010101011010101010101010,
64'b1111111100000000111111110000000001100110011001100110011001100110,
64'b0011001100110011110011001100110001101001100101100110100110010110,
64'b0000000000000000000000000000000011001100001100110011001111001100,
64'b1111000011110000111100001111000000001111000011111111000011110000,
64'b0000000011111111111111110000000000001111111100000000111111110000,
64'b0000000011111111111111110000000011110000111100001111000011110000,
64'b0000000011111111111111110000000011000011001111001100001100111100,
64'b1111111111111111000000000000000011000011001111001100001100111100,
64'b1010101001010101010101011010101011000011110000110011110000111100,
64'b0101010110101010010101011010101001101001011010011001011010010110,
64'b1111000011110000111100001111000010010110100101101001011010010110,
64'b1001011001101001011010011001011010101010010101010101010110101010,
64'b1111111111111111000000000000000001100110011001100110011001100110,
64'b0101010110101010010101011010101010010110100101101001011010010110,
64'b1010010110100101010110100101101010010110011010010110100110010110,
64'b0011110011000011110000110011110000001111000011111111000011110000,
64'b1001100101100110100110010110011001010101101010100101010110101010,
64'b0000000011111111111111110000000010101010010101010101010110101010,
64'b1010101001010101010101011010101011111111000000001111111100000000,
64'b1010101001010101010101011010101011110000000011110000111111110000,
64'b0101010101010101101010101010101011110000000011110000111111110000,
64'b0110011010011001100110010110011000001111111100000000111111110000,
64'b0000111100001111111100001111000001101001100101100110100110010110,
64'b0000111100001111111100001111000001101001100101100110100110010110,
64'b0000111100001111111100001111000000110011001100111100110011001100,
64'b0101010101010101101010101010101010010110100101101001011010010110,
64'b1001100101100110100110010110011011000011001111001100001100111100,
64'b0011001111001100001100111100110000111100110000111100001100111100,
64'b0101101010100101101001010101101001010101101010100101010110101010,
64'b0110100101101001100101101001011010011001100110010110011001100110,
64'b1111111111111111000000000000000000110011001100111100110011001100,
64'b1001100110011001011001100110011001010101010101011010101010101010,
64'b1001100110011001011001100110011000000000111111111111111100000000,
64'b0110011001100110011001100110011010101010010101010101010110101010,
64'b0110100101101001100101101001011010101010010101010101010110101010,
64'b0101010110101010010101011010101000111100110000111100001100111100,
64'b0101010110101010010101011010101000111100110000111100001100111100,
64'b0101010110101010010101011010101011110000111100001111000011110000,
64'b0110011001100110011001100110011001101001100101100110100110010110,
64'b1001011010010110100101101001011000001111111100000000111111110000,
64'b1111000011110000111100001111000001011010101001011010010101011010,
64'b0101101001011010010110100101101010011001100110010110011001100110,
64'b0000111111110000000011111111000000111100001111000011110000111100,
64'b0101010110101010010101011010101001011010010110100101101001011010,
64'b0110100110010110011010011001011001100110011001100110011001100110,
64'b0110100110010110011010011001011001010101010101011010101010101010,
64'b0110100101101001100101101001011010011001100110010110011001100110,
64'b0011110000111100001111000011110010011001100110010110011001100110,
64'b0000111100001111111100001111000001011010101001011010010101011010,
64'b1100001100111100110000110011110001011010101001011010010101011010,
64'b0000000011111111111111110000000001010101101010100101010110101010,
64'b1100001111000011001111000011110000111100110000111100001100111100,
64'b0011110000111100001111000011110011111111000000001111111100000000,
64'b1010101001010101010101011010101011001100001100110011001111001100,
64'b1010010110100101010110100101101010010110100101101001011010010110,
64'b0110011010011001100110010110011010100101010110101010010101011010,
64'b1100110000110011001100111100110000110011110011000011001111001100,
64'b1100001111000011001111000011110000111100001111000011110000111100,
64'b1100001111000011001111000011110011001100110011001100110011001100,
64'b0011110011000011110000110011110010010110100101101001011010010110,
64'b0101101001011010010110100101101010010110100101101001011010010110,
64'b0110100110010110011010011001011001100110100110011001100101100110,
64'b1010101010101010101010101010101001100110100110011001100101100110,
64'b1100110000110011001100111100110010011001100110010110011001100110,
64'b0101101010100101101001010101101011110000000011110000111111110000,
64'b0101101001011010010110100101101010101010101010101010101010101010,
64'b0011001100110011110011001100110011110000111100001111000011110000,
64'b1001100101100110100110010110011011111111111111110000000000000000,
64'b0110100101101001100101101001011010101010010101010101010110101010,
64'b1010010110100101010110100101101011110000000011110000111111110000,
64'b1010010101011010101001010101101011110000111100001111000011110000,
64'b1010010101011010101001010101101000001111111100000000111111110000,
64'b0101101010100101101001010101101000111100110000111100001100111100,
64'b1001100101100110100110010110011000111100001111000011110000111100,
64'b0011110011000011110000110011110001010101010101011010101010101010,
64'b1100110011001100110011001100110010011001011001101001100101100110,
64'b0000111100001111111100001111000010100101010110101010010101011010,
64'b0110011010011001100110010110011001010101101010100101010110101010,
64'b1001100101100110100110010110011010011001011001101001100101100110,
64'b1010010110100101010110100101101010101010010101010101010110101010,
64'b1111111100000000111111110000000010010110011010010110100110010110,
64'b1010010101011010101001010101101011111111111111110000000000000000,
64'b0110011001100110011001100110011001010101010101011010101010101010,
64'b1001100110011001011001100110011010101010101010101010101010101010,
64'b0011001100110011110011001100110011111111111111110000000000000000,
64'b0011001111001100001100111100110000001111111100000000111111110000,
64'b1001011001101001011010011001011001011010010110100101101001011010,
64'b0110011010011001100110010110011001011010010110100101101001011010,
64'b1010101001010101010101011010101010011001011001101001100101100110,
64'b1100110011001100110011001100110011111111111111110000000000000000,
64'b1001011010010110100101101001011011001100110011001100110011001100,
64'b0110100110010110011010011001011011000011001111001100001100111100,
64'b0110011010011001100110010110011010011001100110010110011001100110,
64'b1100001100111100110000110011110010010110011010010110100110010110,
64'b1010101001010101010101011010101010101010101010101010101010101010,
64'b1100001100111100110000110011110001100110011001100110011001100110,
64'b1100001100111100110000110011110001100110011001100110011001100110,
64'b1010010101011010101001010101101000000000000000000000000000000000,
64'b0101101001011010010110100101101010101010010101010101010110101010,
64'b1100001111000011001111000011110000110011110011000011001111001100,
64'b1111111111111111000000000000000000110011110011000011001111001100,
64'b0110100110010110011010011001011011000011110000110011110000111100,
64'b0110100110010110011010011001011000000000000000000000000000000000,
64'b0011110011000011110000110011110001011010010110100101101001011010,
64'b0011110000111100001111000011110000001111111100000000111111110000,
64'b1100001111000011001111000011110010010110100101101001011010010110,
64'b0101101010100101101001010101101010010110011010010110100110010110,
64'b0011001100110011110011001100110001100110011001100110011001100110,
64'b0101101010100101101001010101101000111100001111000011110000111100,
64'b1111000000001111000011111111000000111100001111000011110000111100,
64'b1100110000110011001100111100110000000000000000000000000000000000,
64'b0011001111001100001100111100110000110011001100111100110011001100,
64'b0000111111110000000011111111000010100101101001010101101001011010,
64'b1010101010101010101010101010101000001111000011111111000011110000,
64'b1001011001101001011010011001011000001111111100000000111111110000,
64'b0011110011000011110000110011110010101010101010101010101010101010,
64'b1111000000001111000011111111000000110011110011000011001111001100,
64'b1010010101011010101001010101101011111111000000001111111100000000,
64'b0101101010100101101001010101101010010110011010010110100110010110,
64'b1111000011110000111100001111000010101010101010101010101010101010,
64'b0011110000111100001111000011110011110000111100001111000011110000,
64'b1001100110011001011001100110011011110000111100001111000011110000,
64'b0101010101010101101010101010101011110000111100001111000011110000,
64'b0101101010100101101001010101101011111111000000001111111100000000,
64'b0101101001011010010110100101101000001111000011111111000011110000,
64'b1111111111111111000000000000000001100110011001100110011001100110,
64'b0101101001011010010110100101101011000011001111001100001100111100,
64'b1100110011001100110011001100110001011010010110100101101001011010,
64'b0110100101101001100101101001011011111111000000001111111100000000,
64'b0101010110101010010101011010101011110000111100001111000011110000,
64'b0110011001100110011001100110011011111111000000001111111100000000,
64'b0011001111001100001100111100110010010110011010010110100110010110,
64'b1100001111000011001111000011110001100110011001100110011001100110,
64'b0110100110010110011010011001011011111111000000001111111100000000,
64'b1100001100111100110000110011110011111111000000001111111100000000,
64'b1001100101100110100110010110011011111111000000001111111100000000,
64'b1001100110011001011001100110011011111111111111110000000000000000,
64'b0110011010011001100110010110011011111111000000001111111100000000,
64'b1111111100000000111111110000000010010110100101101001011010010110,
64'b0000111111110000000011111111000011110000000011110000111111110000,
64'b0000000011111111111111110000000000110011110011000011001111001100,
64'b1111000011110000111100001111000011111111111111110000000000000000,
64'b0110011001100110011001100110011011111111000000001111111100000000,
64'b1100001100111100110000110011110000000000000000000000000000000000,
64'b0101101001011010010110100101101010010110011010010110100110010110,
64'b1001100110011001011001100110011010010110100101101001011010010110,
64'b1111000000001111000011111111000011111111111111110000000000000000,
64'b0000111100001111111100001111000011111111111111110000000000000000,
64'b0011110011000011110000110011110011111111111111110000000000000000,
64'b1100001100111100110000110011110000000000000000000000000000000000,
64'b1001011010010110100101101001011001010101010101011010101010101010,
64'b1010101001010101010101011010101011000011001111001100001100111100,
64'b1001011001101001011010011001011000000000111111111111111100000000,
64'b0000111111110000000011111111000010100101101001010101101001011010,
64'b0110011001100110011001100110011000000000000000000000000000000000,
64'b1100001111000011001111000011110001010101010101011010101010101010,
64'b1111000011110000111100001111000000000000000000000000000000000000,
64'b0011001111001100001100111100110000111100110000111100001100111100,
64'b0011110000111100001111000011110001101001100101100110100110010110,
64'b1010101001010101010101011010101000000000000000000000000000000000,
64'b0101010110101010010101011010101010101010101010101010101010101010,
64'b0101101010100101101001010101101010101010101010101010101010101010,
64'b0101101010100101101001010101101010101010101010101010101010101010,
64'b1100001100111100110000110011110011001100110011001100110011001100,
64'b0011001100110011110011001100110001011010101001011010010101011010,
64'b1001011001101001011010011001011011111111111111110000000000000000,
64'b1010101001010101010101011010101010011001011001101001100101100110,
64'b0011110000111100001111000011110010101010101010101010101010101010,
64'b0000111111110000000011111111000011001100110011001100110011001100,
64'b0101010110101010010101011010101010101010101010101010101010101010,
64'b1010010110100101010110100101101011110000000011110000111111110000,
64'b0000111111110000000011111111000010010110011010010110100110010110,
64'b0011001100110011110011001100110000000000000000000000000000000000,
64'b1001100110011001011001100110011011001100110011001100110011001100,
64'b1100110000110011001100111100110011001100110011001100110011001100,
64'b0110011010011001100110010110011011001100110011001100110011001100,
64'b0101101010100101101001010101101011110000111100001111000011110000,
64'b1111000011110000111100001111000011001100001100110011001111001100,
64'b1001011001101001011010011001011010101010101010101010101010101010,
64'b1001100110011001011001100110011001101001011010011001011010010110,
64'b1010010101011010101001010101101011001100110011001100110011001100,
64'b0000000011111111111111110000000011110000111100001111000011110000,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b1001100101100110100110010110011000000000111111111111111100000000,
64'b1010101001010101010101011010101010010110011010010110100110010110,
64'b1111000011110000111100001111000010101010101010101010101010101010,
64'b1001011010010110100101101001011011110000111100001111000011110000,
64'b1010010110100101010110100101101011110000111100001111000011110000,
64'b0110100101101001100101101001011011110000111100001111000011110000,
64'b0110011010011001100110010110011011111111000000001111111100000000,
64'b0101010110101010010101011010101000001111000011111111000011110000,
64'b0011110011000011110000110011110001100110011001100110011001100110,
64'b1001011010010110100101101001011011000011001111001100001100111100,
64'b0110011010011001100110010110011001011010010110100101101001011010,
64'b1111111111111111000000000000000011111111000000001111111100000000,
64'b0101101001011010010110100101101011110000111100001111000011110000,
64'b0000000000000000000000000000000000001111000011111111000011110000,
64'b1001011001101001011010011001011010100101101001010101101001011010,
64'b0000000000000000000000000000000000111100110000111100001100111100,
64'b1010101001010101010101011010101010011001100110010110011001100110,
64'b0101010110101010010101011010101000110011110011000011001111001100,
64'b1001100101100110100110010110011011111111111111110000000000000000,
64'b0000111111110000000011111111000010101010010101010101010110101010,
64'b0110011001100110011001100110011010011001100110010110011001100110,
64'b1111000000001111000011111111000011110000111100001111000011110000,
64'b0101010110101010010101011010101001100110100110011001100101100110,
64'b1100001111000011001111000011110010100101101001010101101001011010,
64'b1111111100000000111111110000000010101010101010101010101010101010,
64'b0011001111001100001100111100110011001100110011001100110011001100,
64'b1010101010101010101010101010101011111111000000001111111100000000,
64'b1010101010101010101010101010101010011001011001101001100101100110,
64'b1010101010101010101010101010101001011010101001011010010101011010,
64'b1001100101100110100110010110011010010110100101101001011010010110,
64'b1100110000110011001100111100110010100101101001010101101001011010,
64'b0101101010100101101001010101101000000000000000000000000000000000,
64'b0000111100001111111100001111000010011001100110010110011001100110,
64'b0101101001011010010110100101101010010110100101101001011010010110,
64'b1111000011110000111100001111000001010101101010100101010110101010,
64'b1100110000110011001100111100110011000011110000110011110000111100,
64'b1100110000110011001100111100110010011001011001101001100101100110,
64'b1010101001010101010101011010101001100110011001100110011001100110,
64'b1100001100111100110000110011110011110000111100001111000011110000,
64'b0110011001100110011001100110011011111111111111110000000000000000,
64'b0101101010100101101001010101101011000011110000110011110000111100,
64'b1100110011001100110011001100110011001100001100110011001111001100,
64'b0110100110010110011010011001011001101001100101100110100110010110,
64'b0101101010100101101001010101101000110011110011000011001111001100,
64'b1111111111111111000000000000000010101010101010101010101010101010,
64'b0101101001011010010110100101101000111100001111000011110000111100,
64'b1111111100000000111111110000000001101001100101100110100110010110,
64'b0000111100001111111100001111000000110011001100111100110011001100,
64'b0101101010100101101001010101101000001111111100000000111111110000,
64'b0110011001100110011001100110011001101001011010011001011010010110,
64'b0110011010011001100110010110011000111100001111000011110000111100,
64'b1001011010010110100101101001011011111111000000001111111100000000,
64'b1001011010010110100101101001011010101010101010101010101010101010,
64'b1100110000110011001100111100110010100101010110101010010101011010,
64'b0101101001011010010110100101101010100101101001010101101001011010,
64'b0011110011000011110000110011110010010110011010010110100110010110,
64'b1100110000110011001100111100110000001111000011111111000011110000,
64'b1010101010101010101010101010101011001100110011001100110011001100,
64'b1001100101100110100110010110011000001111111100000000111111110000,
64'b1111111111111111000000000000000000111100110000111100001100111100,
64'b1111111100000000111111110000000011110000111100001111000011110000,
64'b0110011010011001100110010110011010101010010101010101010110101010,
64'b1001011010010110100101101001011011000011001111001100001100111100,
64'b1100001111000011001111000011110010100101010110101010010101011010,
64'b0110100110010110011010011001011000000000000000000000000000000000,
64'b1100001100111100110000110011110001100110011001100110011001100110,
64'b1001100101100110100110010110011011001100001100110011001111001100,
64'b1001100101100110100110010110011000110011110011000011001111001100,
64'b0101101001011010010110100101101010010110011010010110100110010110,
64'b1111000000001111000011111111000001010101101010100101010110101010,
64'b1111111100000000111111110000000001011010010110100101101001011010,
64'b1100110000110011001100111100110000000000111111111111111100000000,
64'b0110011001100110011001100110011011110000000011110000111111110000,
64'b1010010101011010101001010101101001010101101010100101010110101010,
64'b1001011001101001011010011001011000110011001100111100110011001100,
64'b1010101001010101010101011010101001011010101001011010010101011010,
64'b1111000011110000111100001111000011001100001100110011001111001100,
64'b0101101001011010010110100101101000000000000000000000000000000000,
64'b1111000000001111000011111111000010010110100101101001011010010110,
64'b0101010110101010010101011010101000001111000011111111000011110000,
64'b1100001111000011001111000011110010100101101001010101101001011010,
64'b1001100110011001011001100110011000111100110000111100001100111100,
64'b0101010101010101101010101010101010011001100110010110011001100110,
64'b1100110000110011001100111100110000110011110011000011001111001100,
64'b0000000011111111111111110000000011111111111111110000000000000000,
64'b1111000011110000111100001111000010101010010101010101010110101010,
64'b0011110000111100001111000011110010011001100110010110011001100110,
64'b0110100101101001100101101001011011110000111100001111000011110000,
64'b0101101001011010010110100101101001100110100110011001100101100110,
64'b1010101010101010101010101010101010100101101001010101101001011010,
64'b0000000000000000000000000000000010101010101010101010101010101010,
64'b0000000011111111111111110000000011000011001111001100001100111100,
64'b1001100110011001011001100110011001101001011010011001011010010110,
64'b0000111111110000000011111111000010011001011001101001100101100110,
64'b1001011010010110100101101001011011110000111100001111000011110000,
64'b0110011001100110011001100110011011000011001111001100001100111100,
64'b1010010110100101010110100101101000111100110000111100001100111100,
64'b0101010101010101101010101010101000001111111100000000111111110000,
64'b0101010110101010010101011010101011111111111111110000000000000000,
64'b0000111111110000000011111111000001100110100110011001100101100110,
64'b1100001100111100110000110011110000000000000000000000000000000000,
64'b1001100101100110100110010110011000000000000000000000000000000000,
64'b1100110011001100110011001100110001100110011001100110011001100110,
64'b0000000000000000000000000000000001010101101010100101010110101010,
64'b0101010101010101101010101010101001011010101001011010010101011010,
64'b0000000011111111111111110000000001010101010101011010101010101010,
64'b1010101001010101010101011010101001101001011010011001011010010110,
64'b0110100101101001100101101001011001010101010101011010101010101010,
64'b0110100110010110011010011001011010100101101001010101101001011010,
64'b1010101010101010101010101010101001101001011010011001011010010110,
64'b0110100110010110011010011001011010100101101001010101101001011010,
64'b1111111111111111000000000000000001100110011001100110011001100110,
64'b1111000011110000111100001111000010011001011001101001100101100110,
64'b1010010110100101010110100101101011111111000000001111111100000000,
64'b0000000000000000000000000000000011000011110000110011110000111100,
64'b0000111111110000000011111111000011000011001111001100001100111100,
64'b0011001111001100001100111100110011111111000000001111111100000000,
64'b0110011001100110011001100110011001100110100110011001100101100110,
64'b1100001100111100110000110011110001100110011001100110011001100110,
64'b1001100110011001011001100110011001101001100101100110100110010110,
64'b1100001111000011001111000011110001100110011001100110011001100110,
64'b1100001111000011001111000011110010011001011001101001100101100110,
64'b0101010110101010010101011010101001101001100101100110100110010110,
64'b0011001100110011110011001100110010011001011001101001100101100110,
64'b0110011001100110011001100110011010010110100101101001011010010110,
64'b1010010110100101010110100101101011000011110000110011110000111100,
64'b0110011001100110011001100110011011111111111111110000000000000000,
64'b0110100101101001100101101001011000001111111100000000111111110000,
64'b1111111111111111000000000000000001011010101001011010010101011010,
64'b1100001100111100110000110011110000000000000000000000000000000000,
64'b0011110000111100001111000011110001101001011010011001011010010110,
64'b1111000000001111000011111111000010010110100101101001011010010110,
64'b0011110000111100001111000011110000111100110000111100001100111100,
64'b1010010101011010101001010101101000111100001111000011110000111100,
64'b1010010101011010101001010101101011000011110000110011110000111100,
64'b1001100110011001011001100110011000111100110000111100001100111100,
64'b1111000011110000111100001111000011000011110000110011110000111100,
64'b1001011010010110100101101001011011000011001111001100001100111100,
64'b0011001111001100001100111100110000001111111100000000111111110000,
64'b1001011010010110100101101001011010101010101010101010101010101010,
64'b1100001100111100110000110011110010101010010101010101010110101010,
64'b1010101010101010101010101010101011001100001100110011001111001100,
64'b1010010101011010101001010101101010101010101010101010101010101010,
64'b1010010101011010101001010101101001101001100101100110100110010110,
64'b1001011010010110100101101001011011111111111111110000000000000000,
64'b1010010101011010101001010101101011110000000011110000111111110000,
64'b0110011001100110011001100110011000001111000011111111000011110000,
64'b1001100110011001011001100110011001011010010110100101101001011010,
64'b1010010101011010101001010101101011000011110000110011110000111100,
64'b0101101001011010010110100101101010101010101010101010101010101010,
64'b1010010101011010101001010101101000111100110000111100001100111100,
64'b1111111100000000111111110000000011110000111100001111000011110000,
64'b1001011010010110100101101001011010011001011001101001100101100110,
64'b0011001111001100001100111100110011110000111100001111000011110000,
64'b0011001111001100001100111100110001011010101001011010010101011010,
64'b0000000000000000000000000000000001010101101010100101010110101010,
64'b1100110000110011001100111100110010010110011010010110100110010110,
64'b0101010101010101101010101010101000000000000000000000000000000000,
64'b1100110000110011001100111100110010101010010101010101010110101010,
64'b1001011001101001011010011001011001010101101010100101010110101010,
64'b0110100110010110011010011001011010011001011001101001100101100110,
64'b1111111111111111000000000000000000001111111100000000111111110000,
64'b0011110000111100001111000011110001100110011001100110011001100110,
64'b1010101001010101010101011010101011110000000011110000111111110000,
64'b0000111111110000000011111111000001010101101010100101010110101010,
64'b1001011010010110100101101001011011000011110000110011110000111100,
64'b1100110011001100110011001100110011111111000000001111111100000000,
64'b1111000000001111000011111111000011001100001100110011001111001100,
64'b0011001111001100001100111100110001100110011001100110011001100110,
64'b1010010110100101010110100101101000111100110000111100001100111100,
64'b1111000000001111000011111111000010101010101010101010101010101010,
64'b1010010110100101010110100101101000110011001100111100110011001100,
64'b0011110000111100001111000011110010011001100110010110011001100110,
64'b1100001111000011001111000011110011000011110000110011110000111100,
64'b1001100101100110100110010110011000000000111111111111111100000000,
64'b1010101010101010101010101010101000111100001111000011110000111100,
64'b0101010101010101101010101010101000000000111111111111111100000000,
64'b0101101001011010010110100101101010011001100110010110011001100110,
64'b1001011010010110100101101001011000001111111100000000111111110000,
64'b0011001100110011110011001100110001010101010101011010101010101010,
64'b1111111111111111000000000000000000001111000011111111000011110000,
64'b0110100110010110011010011001011010010110100101101001011010010110,
64'b0011001111001100001100111100110011110000000011110000111111110000,
64'b1010101001010101010101011010101001100110011001100110011001100110,
64'b1001100101100110100110010110011011110000111100001111000011110000,
64'b1010010101011010101001010101101010010110100101101001011010010110,
64'b0000111111110000000011111111000010100101010110101010010101011010,
64'b0110100101101001100101101001011001010101010101011010101010101010,
64'b1100110011001100110011001100110010100101010110101010010101011010,
64'b1100110011001100110011001100110011111111111111110000000000000000,
64'b1001100101100110100110010110011010010110100101101001011010010110,
64'b1100001100111100110000110011110010101010010101010101010110101010,
64'b1111000011110000111100001111000011001100110011001100110011001100,
64'b1010101010101010101010101010101001010101101010100101010110101010,
64'b0110100110010110011010011001011001101001100101100110100110010110,
64'b1010010110100101010110100101101000000000111111111111111100000000,
64'b0011001100110011110011001100110010010110100101101001011010010110,
64'b0110100101101001100101101001011011111111000000001111111100000000,
64'b1100110000110011001100111100110011000011001111001100001100111100,
64'b0000000011111111111111110000000011001100001100110011001111001100,
64'b1100001100111100110000110011110011001100110011001100110011001100,
64'b0101101001011010010110100101101001100110100110011001100101100110,
64'b1111000011110000111100001111000000000000000000000000000000000000,
64'b1100001111000011001111000011110001101001100101100110100110010110,
64'b1111000000001111000011111111000000110011001100111100110011001100,
64'b1111111100000000111111110000000001011010010110100101101001011010,
64'b1100110011001100110011001100110000110011001100111100110011001100,
64'b1100001100111100110000110011110011000011001111001100001100111100,
64'b0011001111001100001100111100110011111111111111110000000000000000,
64'b0101101001011010010110100101101001101001100101100110100110010110,
64'b0110100110010110011010011001011011111111111111110000000000000000,
64'b1010010110100101010110100101101011110000000011110000111111110000,
64'b0101010101010101101010101010101000001111000011111111000011110000,
64'b0101101010100101101001010101101001011010010110100101101001011010,
64'b0011001111001100001100111100110011000011110000110011110000111100,
64'b1111111100000000111111110000000010101010101010101010101010101010,
64'b0000111111110000000011111111000000111100110000111100001100111100,
64'b1010101001010101010101011010101011110000111100001111000011110000,
64'b0101010101010101101010101010101010011001011001101001100101100110,
64'b1111000011110000111100001111000011110000111100001111000011110000,
64'b0000111111110000000011111111000010100101010110101010010101011010,
64'b1001011010010110100101101001011011111111000000001111111100000000,
64'b1001011010010110100101101001011001100110100110011001100101100110,
64'b0011001100110011110011001100110011110000111100001111000011110000,
64'b1111111111111111000000000000000000001111000011111111000011110000,
64'b0000111111110000000011111111000000111100110000111100001100111100,
64'b1111111100000000111111110000000010011001011001101001100101100110,
64'b0011001100110011110011001100110010101010010101010101010110101010,
64'b1010010110100101010110100101101011000011001111001100001100111100,
64'b0110100101101001100101101001011001101001011010011001011010010110,
64'b0011001100110011110011001100110000001111000011111111000011110000,
64'b1111000011110000111100001111000001010101010101011010101010101010,
64'b1111000000001111000011111111000011001100110011001100110011001100,
64'b1001011010010110100101101001011010011001011001101001100101100110,
64'b1111111100000000111111110000000011111111111111110000000000000000,
64'b0101010110101010010101011010101011000011110000110011110000111100,
64'b1100001111000011001111000011110001010101101010100101010110101010,
64'b0101010101010101101010101010101011111111000000001111111100000000,
64'b1010010110100101010110100101101001011010101001011010010101011010,
64'b0000000011111111111111110000000001101001011010011001011010010110,
64'b1100001111000011001111000011110000110011001100111100110011001100,
64'b0011110011000011110000110011110001011010101001011010010101011010,
64'b0000000011111111111111110000000011000011001111001100001100111100,
64'b0110100101101001100101101001011001010101101010100101010110101010,
64'b1010010101011010101001010101101001100110011001100110011001100110,
64'b1111000011110000111100001111000001011010010110100101101001011010,
64'b1111111100000000111111110000000000111100001111000011110000111100,
64'b1100001111000011001111000011110000000000000000000000000000000000,
64'b1010010110100101010110100101101010100101010110101010010101011010,
64'b0011110011000011110000110011110010011001100110010110011001100110,
64'b1001100110011001011001100110011011111111111111110000000000000000,
64'b1001011010010110100101101001011011001100001100110011001111001100,
64'b1010101001010101010101011010101001101001100101100110100110010110,
64'b1001011001101001011010011001011001011010010110100101101001011010,
64'b1111111100000000111111110000000001100110100110011001100101100110,
64'b0011110000111100001111000011110001011010101001011010010101011010,
64'b0101101010100101101001010101101000110011001100111100110011001100,
64'b1001011001101001011010011001011000111100001111000011110000111100,
64'b0000111100001111111100001111000000110011110011000011001111001100,
64'b1001011010010110100101101001011000001111111100000000111111110000,
64'b0000111111110000000011111111000010101010101010101010101010101010,
64'b1001100101100110100110010110011011001100001100110011001111001100,
64'b0101101010100101101001010101101000111100001111000011110000111100,
64'b1001011010010110100101101001011010101010101010101010101010101010,
64'b0110100110010110011010011001011010100101101001010101101001011010,
64'b0011001100110011110011001100110010010110011010010110100110010110,
64'b1001011001101001011010011001011000110011110011000011001111001100,
64'b0101010101010101101010101010101011000011110000110011110000111100,
64'b0000111111110000000011111111000001100110100110011001100101100110,
64'b1100110000110011001100111100110001011010010110100101101001011010,
64'b1001011001101001011010011001011010100101010110101010010101011010,
64'b0101010110101010010101011010101000001111000011111111000011110000,
64'b0110100110010110011010011001011011111111000000001111111100000000,
64'b0011110011000011110000110011110011001100110011001100110011001100,
64'b0101010101010101101010101010101000001111000011111111000011110000,
64'b1111111100000000111111110000000010100101010110101010010101011010,
64'b1001011001101001011010011001011011001100110011001100110011001100,
64'b0011001100110011110011001100110000110011110011000011001111001100,
64'b0000111111110000000011111111000010010110011010010110100110010110,
64'b1010010101011010101001010101101010100101101001010101101001011010,
64'b1100001111000011001111000011110000001111111100000000111111110000,
64'b1100001100111100110000110011110001101001011010011001011010010110,
64'b0011110000111100001111000011110010011001011001101001100101100110,
64'b0110011010011001100110010110011011001100001100110011001111001100,
64'b0110100110010110011010011001011011111111000000001111111100000000,
64'b0101010110101010010101011010101010101010101010101010101010101010,
64'b0110011010011001100110010110011011110000111100001111000011110000,
64'b1111000011110000111100001111000011111111000000001111111100000000,
64'b0110011001100110011001100110011001100110100110011001100101100110,
64'b1100001100111100110000110011110011110000111100001111000011110000,
64'b0101010110101010010101011010101000001111000011111111000011110000,
64'b0101010101010101101010101010101000111100110000111100001100111100,
64'b1111111100000000111111110000000010011001011001101001100101100110,
64'b1010101001010101010101011010101010101010010101010101010110101010,
64'b0011001111001100001100111100110011000011001111001100001100111100,
64'b0011110011000011110000110011110001101001011010011001011010010110,
64'b0011001100110011110011001100110000001111000011111111000011110000,
64'b0110011001100110011001100110011001010101010101011010101010101010,
64'b0101101001011010010110100101101011001100110011001100110011001100,
64'b1100001111000011001111000011110001101001100101100110100110010110,
64'b0101010110101010010101011010101001101001011010011001011010010110,
64'b0011110000111100001111000011110011110000111100001111000011110000,
64'b1111000000001111000011111111000010101010010101010101010110101010,
64'b0011001100110011110011001100110011110000111100001111000011110000,
64'b1100110011001100110011001100110010100101101001010101101001011010,
64'b0101010101010101101010101010101001011010010110100101101001011010,
64'b0011001100110011110011001100110010010110100101101001011010010110,
64'b1010010110100101010110100101101000110011110011000011001111001100,
64'b1111000000001111000011111111000011110000000011110000111111110000,
64'b0101101001011010010110100101101010100101010110101010010101011010,
64'b1001011010010110100101101001011010010110011010010110100110010110,
64'b0011001111001100001100111100110011001100110011001100110011001100,
64'b1001100101100110100110010110011000000000111111111111111100000000,
64'b0000111100001111111100001111000001010101101010100101010110101010,
64'b0011110011000011110000110011110001100110100110011001100101100110,
64'b1111111100000000111111110000000011001100110011001100110011001100,
64'b0101010110101010010101011010101001011010010110100101101001011010,
64'b1010010101011010101001010101101011001100110011001100110011001100,
64'b1111111111111111000000000000000010101010010101010101010110101010,
64'b1111111111111111000000000000000001100110100110011001100101100110,
64'b1111000000001111000011111111000001100110011001100110011001100110,
64'b1001100101100110100110010110011000110011110011000011001111001100,
64'b0110100110010110011010011001011010010110011010010110100110010110,
64'b0011001100110011110011001100110011001100110011001100110011001100,
64'b0110011001100110011001100110011011001100110011001100110011001100,
64'b1111111111111111000000000000000001010101010101011010101010101010,
64'b0110100110010110011010011001011010011001100110010110011001100110,
64'b0110100110010110011010011001011011000011110000110011110000111100,
64'b1010101010101010101010101010101001011010010110100101101001011010,
64'b0011110011000011110000110011110000110011110011000011001111001100,
64'b0011001100110011110011001100110011110000111100001111000011110000,
64'b0011001100110011110011001100110000110011001100111100110011001100,
64'b0000111100001111111100001111000001101001011010011001011010010110,
64'b1100001100111100110000110011110010010110100101101001011010010110,
64'b0101101001011010010110100101101000001111000011111111000011110000,
64'b1100110000110011001100111100110000111100110000111100001100111100,
64'b0000000011111111111111110000000001011010010110100101101001011010,
64'b0000000000000000000000000000000011110000111100001111000011110000,
64'b1010101010101010101010101010101011001100110011001100110011001100,
64'b1001011001101001011010011001011010010110100101101001011010010110,
64'b0011110011000011110000110011110010100101010110101010010101011010,
64'b1100110011001100110011001100110010011001011001101001100101100110,
64'b1111000000001111000011111111000000001111000011111111000011110000,
64'b0101101001011010010110100101101011111111000000001111111100000000,
64'b0101101001011010010110100101101011110000111100001111000011110000,
64'b0101010110101010010101011010101001101001100101100110100110010110,
64'b0101101010100101101001010101101001101001100101100110100110010110,
64'b0011001111001100001100111100110011111111000000001111111100000000,
64'b0000111100001111111100001111000001011010101001011010010101011010,
64'b0101010101010101101010101010101010011001011001101001100101100110,
64'b1010101010101010101010101010101011111111000000001111111100000000,
64'b1111000011110000111100001111000001100110011001100110011001100110,
64'b1010101001010101010101011010101001010101101010100101010110101010,
64'b0110100110010110011010011001011011111111000000001111111100000000,
64'b1010010110100101010110100101101000111100001111000011110000111100,
64'b0000111100001111111100001111000011110000111100001111000011110000,
64'b0110011001100110011001100110011010101010010101010101010110101010,
64'b0000000011111111111111110000000011001100001100110011001111001100,
64'b1001011010010110100101101001011010011001011001101001100101100110,
64'b1010010101011010101001010101101001010101101010100101010110101010,
64'b1001011010010110100101101001011011001100110011001100110011001100,
64'b0000111111110000000011111111000000111100110000111100001100111100,
64'b1001011001101001011010011001011010011001011001101001100101100110,
64'b1111000011110000111100001111000010010110100101101001011010010110,
64'b0110100110010110011010011001011010010110100101101001011010010110,
64'b1010010110100101010110100101101000110011001100111100110011001100,
64'b1010010101011010101001010101101011111111111111110000000000000000,
64'b1100110000110011001100111100110000001111111100000000111111110000,
64'b0101101001011010010110100101101011111111000000001111111100000000,
64'b0110100110010110011010011001011000110011001100111100110011001100,
64'b1100110011001100110011001100110010100101101001010101101001011010,
64'b1100110000110011001100111100110001101001011010011001011010010110,
64'b1010010101011010101001010101101000110011001100111100110011001100,
64'b1111000000001111000011111111000011110000111100001111000011110000,
64'b1111000000001111000011111111000011110000000011110000111111110000,
64'b1100110011001100110011001100110001101001011010011001011010010110,
64'b1100001100111100110000110011110011000011001111001100001100111100,
64'b0000000011111111111111110000000011000011001111001100001100111100,
64'b1010010101011010101001010101101011110000111100001111000011110000,
64'b0101010110101010010101011010101010101010101010101010101010101010,
64'b1111000011110000111100001111000010101010010101010101010110101010,
64'b1001011010010110100101101001011011111111111111110000000000000000,
64'b1100001111000011001111000011110011110000111100001111000011110000,
64'b1100001111000011001111000011110010011001011001101001100101100110,
64'b1010101010101010101010101010101001101001100101100110100110010110,
64'b0000111111110000000011111111000001011010010110100101101001011010,
64'b0011001111001100001100111100110001010101101010100101010110101010,
64'b0101101010100101101001010101101000000000111111111111111100000000,
64'b1010101001010101010101011010101001101001100101100110100110010110,
64'b1001100101100110100110010110011010100101010110101010010101011010,
64'b0101010101010101101010101010101011110000000011110000111111110000,
64'b0110011010011001100110010110011011111111000000001111111100000000,
64'b0011001100110011110011001100110011001100110011001100110011001100,
64'b1111111100000000111111110000000000110011001100111100110011001100,
64'b1100001100111100110000110011110010101010101010101010101010101010,
64'b0000111111110000000011111111000001010101101010100101010110101010,
64'b1010010101011010101001010101101011000011110000110011110000111100,
64'b0110011001100110011001100110011000111100110000111100001100111100,
64'b0000000011111111111111110000000000110011110011000011001111001100,
64'b0000111100001111111100001111000000110011001100111100110011001100,
64'b1100110000110011001100111100110011111111111111110000000000000000,
64'b1001100110011001011001100110011010010110011010010110100110010110,
64'b1001011010010110100101101001011000110011110011000011001111001100,
64'b0110011001100110011001100110011010101010010101010101010110101010,
64'b0110100101101001100101101001011001010101010101011010101010101010,
64'b0101101001011010010110100101101011110000111100001111000011110000,
64'b0101010101010101101010101010101011110000111100001111000011110000,
64'b1111000000001111000011111111000001100110011001100110011001100110,
64'b0000000011111111111111110000000000110011001100111100110011001100,
64'b1100110000110011001100111100110000001111111100000000111111110000,
64'b0011110000111100001111000011110001011010101001011010010101011010,
64'b1111111111111111000000000000000010100101101001010101101001011010,
64'b0101010110101010010101011010101011110000111100001111000011110000,
64'b1010010110100101010110100101101010101010101010101010101010101010,
64'b1001011010010110100101101001011010010110011010010110100110010110,
64'b0110100110010110011010011001011001011010010110100101101001011010,
64'b1001011010010110100101101001011010011001100110010110011001100110,
64'b1100001100111100110000110011110001100110011001100110011001100110,
64'b1001100101100110100110010110011001010101101010100101010110101010,
64'b1100110011001100110011001100110011111111000000001111111100000000,
64'b1010101001010101010101011010101000111100001111000011110000111100,
64'b0101010101010101101010101010101011110000111100001111000011110000,
64'b1010010110100101010110100101101010101010010101010101010110101010,
64'b1010010101011010101001010101101011001100001100110011001111001100,
64'b0000000000000000000000000000000010011001011001101001100101100110,
64'b1001100110011001011001100110011001010101101010100101010110101010,
64'b0011001111001100001100111100110011001100110011001100110011001100,
64'b0110100110010110011010011001011000111100110000111100001100111100,
64'b1100001100111100110000110011110010011001011001101001100101100110,
64'b0101101010100101101001010101101011000011110000110011110000111100,
64'b1111111100000000111111110000000001010101101010100101010110101010,
64'b1100001100111100110000110011110000110011001100111100110011001100,
64'b0101101010100101101001010101101010100101101001010101101001011010,
64'b1111111111111111000000000000000001011010101001011010010101011010,
64'b1100001111000011001111000011110000001111111100000000111111110000,
64'b0011110011000011110000110011110010101010010101010101010110101010,
64'b0110011010011001100110010110011001101001011010011001011010010110,
64'b0110100110010110011010011001011001010101101010100101010110101010,
64'b1001100101100110100110010110011010011001011001101001100101100110,
64'b1010101010101010101010101010101000001111000011111111000011110000,
64'b0110100110010110011010011001011010010110011010010110100110010110,
64'b0101010110101010010101011010101011111111000000001111111100000000,
64'b1001011010010110100101101001011010100101010110101010010101011010,
64'b1010101001010101010101011010101010011001100110010110011001100110,
64'b0011001100110011110011001100110011110000111100001111000011110000,
64'b1001011010010110100101101001011010011001011001101001100101100110,
64'b0101010101010101101010101010101001100110100110011001100101100110,
64'b0110011010011001100110010110011010101010010101010101010110101010,
64'b0110011001100110011001100110011000110011001100111100110011001100,
64'b0000111111110000000011111111000001101001100101100110100110010110,
64'b1111111111111111000000000000000010011001100110010110011001100110,
64'b0101101010100101101001010101101011000011110000110011110000111100,
64'b0110011001100110011001100110011011111111000000001111111100000000,
64'b0101010101010101101010101010101010010110011010010110100110010110,
64'b1001100101100110100110010110011010101010101010101010101010101010,
64'b0011001100110011110011001100110011001100001100110011001111001100,
64'b1100110000110011001100111100110000111100001111000011110000111100,
64'b1001100101100110100110010110011001010101101010100101010110101010,
64'b0011001100110011110011001100110011000011110000110011110000111100,
64'b0011001100110011110011001100110011000011110000110011110000111100,
64'b1010101010101010101010101010101010011001100110010110011001100110,
64'b1010101001010101010101011010101001011010010110100101101001011010,
64'b0110011001100110011001100110011010010110011010010110100110010110,
64'b0110100110010110011010011001011000111100001111000011110000111100,
64'b1111111111111111000000000000000010100101010110101010010101011010,
64'b0011110000111100001111000011110001010101010101011010101010101010,
64'b1010010101011010101001010101101000111100110000111100001100111100,
64'b1100001100111100110000110011110001100110011001100110011001100110,
64'b1111000011110000111100001111000010100101101001010101101001011010,
64'b1010010110100101010110100101101010100101010110101010010101011010,
64'b0110100101101001100101101001011000110011001100111100110011001100,
64'b1111000011110000111100001111000000001111111100000000111111110000,
64'b0101101001011010010110100101101010100101010110101010010101011010,
64'b0110011001100110011001100110011010010110100101101001011010010110,
64'b0011001100110011110011001100110010011001011001101001100101100110,
64'b1001011010010110100101101001011000111100110000111100001100111100,
64'b0011110011000011110000110011110010100101010110101010010101011010,
64'b0000000000000000000000000000000011001100001100110011001111001100,
64'b1010010101011010101001010101101011001100110011001100110011001100,
64'b1100110000110011001100111100110001011010101001011010010101011010,
64'b0000111111110000000011111111000010010110100101101001011010010110,
64'b0000111100001111111100001111000010011001011001101001100101100110,
64'b1100110011001100110011001100110001100110100110011001100101100110,
64'b1010101010101010101010101010101011110000111100001111000011110000,
64'b0000111100001111111100001111000010101010010101010101010110101010,
64'b1100110000110011001100111100110011001100001100110011001111001100,
64'b1111111111111111000000000000000011000011001111001100001100111100,
64'b1100110000110011001100111100110011000011110000110011110000111100,
64'b0000111100001111111100001111000011110000000011110000111111110000,
64'b1001100110011001011001100110011001100110100110011001100101100110,
64'b0011001111001100001100111100110000001111000011111111000011110000,
64'b0110011010011001100110010110011001011010010110100101101001011010,
64'b0110011010011001100110010110011011001100001100110011001111001100,
64'b0000000000000000000000000000000001101001100101100110100110010110,
64'b0000111100001111111100001111000011000011110000110011110000111100,
64'b1010010101011010101001010101101011000011110000110011110000111100,
64'b0000111111110000000011111111000001010101101010100101010110101010,
64'b1010010110100101010110100101101000110011001100111100110011001100,
64'b0101101001011010010110100101101010100101101001010101101001011010,
64'b0110100101101001100101101001011001011010101001011010010101011010,
64'b1001100101100110100110010110011000001111111100000000111111110000,
64'b0011001100110011110011001100110010101010010101010101010110101010,
64'b1111111100000000111111110000000001101001011010011001011010010110,
64'b0011110011000011110000110011110001010101101010100101010110101010,
64'b0110100101101001100101101001011010011001011001101001100101100110,
64'b0000000011111111111111110000000000001111000011111111000011110000,
64'b1111111100000000111111110000000001101001100101100110100110010110,
64'b1111111100000000111111110000000001010101010101011010101010101010,
64'b0110011010011001100110010110011001011010010110100101101001011010,
64'b0000000011111111111111110000000001011010101001011010010101011010,
64'b0011001111001100001100111100110010101010010101010101010110101010,
64'b1001100101100110100110010110011001100110100110011001100101100110,
64'b1100001100111100110000110011110010100101010110101010010101011010,
64'b0110100101101001100101101001011010010110100101101001011010010110,
64'b1111000011110000111100001111000001010101101010100101010110101010,
64'b0101010101010101101010101010101000000000000000000000000000000000,
64'b1111000000001111000011111111000000000000111111111111111100000000,
64'b0110100110010110011010011001011001101001011010011001011010010110,
64'b0101010101010101101010101010101010010110100101101001011010010110,
64'b1010101010101010101010101010101000111100001111000011110000111100,
64'b0000111111110000000011111111000010010110011010010110100110010110,
64'b0011110011000011110000110011110001100110011001100110011001100110,
64'b1001011001101001011010011001011000001111000011111111000011110000,
64'b1111111100000000111111110000000011000011001111001100001100111100,
64'b0011110000111100001111000011110010010110100101101001011010010110,
64'b0011001111001100001100111100110010100101010110101010010101011010,
64'b1111111111111111000000000000000011111111111111110000000000000000,
64'b0011001100110011110011001100110001010101101010100101010110101010,
64'b1010010101011010101001010101101001101001100101100110100110010110,
64'b0011001100110011110011001100110001100110100110011001100101100110,
64'b0011110011000011110000110011110011000011001111001100001100111100,
64'b1010010101011010101001010101101000000000000000000000000000000000,
64'b0011001111001100001100111100110001011010010110100101101001011010,
64'b0101101001011010010110100101101000111100110000111100001100111100,
64'b0000111100001111111100001111000010010110100101101001011010010110,
64'b0101010101010101101010101010101011111111000000001111111100000000,
64'b0000111111110000000011111111000001011010101001011010010101011010,
64'b1111000000001111000011111111000011000011001111001100001100111100,
64'b1100110011001100110011001100110011001100001100110011001111001100,
64'b0011110011000011110000110011110000000000000000000000000000000000,
64'b0011110011000011110000110011110010011001100110010110011001100110,
64'b0000111100001111111100001111000000111100110000111100001100111100,
64'b0110100110010110011010011001011011000011110000110011110000111100,
64'b1111000000001111000011111111000001011010101001011010010101011010,
64'b0000111100001111111100001111000000000000000000000000000000000000,
64'b1010010101011010101001010101101000110011110011000011001111001100,
64'b0011001111001100001100111100110011110000000011110000111111110000,
64'b1111111100000000111111110000000001101001100101100110100110010110,
64'b0110011001100110011001100110011011111111111111110000000000000000,
64'b1010101001010101010101011010101011001100001100110011001111001100,
64'b0000000011111111111111110000000001011010101001011010010101011010,
64'b0101101001011010010110100101101000001111000011111111000011110000,
64'b1111000000001111000011111111000010101010101010101010101010101010,
64'b0101101010100101101001010101101000111100001111000011110000111100,
64'b0101010110101010010101011010101001011010101001011010010101011010,
64'b1001011001101001011010011001011010100101010110101010010101011010,
64'b0000000011111111111111110000000001100110100110011001100101100110,
64'b0101010110101010010101011010101010101010101010101010101010101010,
64'b1001100101100110100110010110011011110000111100001111000011110000,
64'b0101010110101010010101011010101011110000111100001111000011110000,
64'b0000000011111111111111110000000001101001011010011001011010010110,
64'b1111111100000000111111110000000011000011001111001100001100111100,
64'b0110100110010110011010011001011011111111000000001111111100000000,
64'b1010101010101010101010101010101010011001011001101001100101100110,
64'b0101101010100101101001010101101010010110011010010110100110010110,
64'b0011110000111100001111000011110001011010101001011010010101011010,
64'b0000000000000000000000000000000001101001011010011001011010010110,
64'b1111000000001111000011111111000010100101101001010101101001011010,
64'b1010010110100101010110100101101011111111111111110000000000000000,
64'b1111111111111111000000000000000001101001011010011001011010010110,
64'b1111000000001111000011111111000000001111111100000000111111110000,
64'b0110100110010110011010011001011010101010101010101010101010101010,
64'b0110100110010110011010011001011011111111000000001111111100000000,
64'b0000000011111111111111110000000011000011001111001100001100111100,
64'b1001011001101001011010011001011001011010101001011010010101011010,
64'b0110011001100110011001100110011011111111111111110000000000000000,
64'b0011001100110011110011001100110011000011110000110011110000111100,
64'b0000111111110000000011111111000000111100110000111100001100111100,
64'b1001100110011001011001100110011001100110100110011001100101100110,
64'b0110011010011001100110010110011001101001100101100110100110010110,
64'b0110100101101001100101101001011010011001011001101001100101100110,
64'b0000000000000000000000000000000010101010101010101010101010101010,
64'b0000000000000000000000000000000001101001100101100110100110010110,
64'b1100001111000011001111000011110010101010010101010101010110101010,
64'b0011110000111100001111000011110011001100110011001100110011001100,
64'b1100110011001100110011001100110001010101010101011010101010101010,
64'b0000000011111111111111110000000011110000000011110000111111110000,
64'b0101010101010101101010101010101011001100001100110011001111001100,
64'b1100110000110011001100111100110010101010101010101010101010101010,
64'b0000111100001111111100001111000010100101010110101010010101011010,
64'b0110100110010110011010011001011001011010101001011010010101011010,
64'b0000000011111111111111110000000001101001011010011001011010010110,
64'b0000111111110000000011111111000010010110011010010110100110010110,
64'b0000000000000000000000000000000011000011110000110011110000111100,
64'b0011001111001100001100111100110011001100110011001100110011001100,
64'b1010101010101010101010101010101000111100110000111100001100111100,
64'b0110011001100110011001100110011000110011001100111100110011001100,
64'b1111000011110000111100001111000001011010010110100101101001011010,
64'b0101101001011010010110100101101001100110011001100110011001100110,
64'b1111111111111111000000000000000010101010010101010101010110101010,
64'b0110011001100110011001100110011010100101101001010101101001011010,
64'b1010010110100101010110100101101001100110011001100110011001100110,
64'b0101010110101010010101011010101011001100001100110011001111001100,
64'b1001011001101001011010011001011011001100001100110011001111001100,
64'b1111111111111111000000000000000001101001100101100110100110010110,
64'b1010101001010101010101011010101010010110011010010110100110010110,
64'b0000000000000000000000000000000010100101010110101010010101011010,
64'b0000111100001111111100001111000001011010010110100101101001011010,
64'b1100110011001100110011001100110011110000000011110000111111110000,
64'b0011110000111100001111000011110001011010010110100101101001011010,
64'b1111111100000000111111110000000010011001011001101001100101100110,
64'b0011001111001100001100111100110010010110100101101001011010010110,
64'b0000000000000000000000000000000000110011001100111100110011001100,
64'b1001011010010110100101101001011010011001011001101001100101100110,
64'b0011001111001100001100111100110010010110100101101001011010010110,
64'b1001100110011001011001100110011000001111000011111111000011110000,
64'b0011110011000011110000110011110010100101101001010101101001011010,
64'b1010101010101010101010101010101010010110011010010110100110010110,
64'b1001100110011001011001100110011000111100110000111100001100111100,
64'b1010101010101010101010101010101001100110100110011001100101100110,
64'b1111111100000000111111110000000000110011110011000011001111001100,
64'b0101101001011010010110100101101000000000111111111111111100000000,
64'b0000111111110000000011111111000010011001011001101001100101100110,
64'b0000000000000000000000000000000000111100001111000011110000111100,
64'b1010010110100101010110100101101011000011001111001100001100111100,
64'b0000000000000000000000000000000011110000111100001111000011110000,
64'b1100001100111100110000110011110001101001011010011001011010010110,
64'b0000111100001111111100001111000011000011001111001100001100111100,
64'b0011110000111100001111000011110011111111000000001111111100000000,
64'b0101101010100101101001010101101010011001011001101001100101100110,
64'b0110011001100110011001100110011010010110011010010110100110010110,
64'b0011110000111100001111000011110001011010101001011010010101011010,
64'b0110011001100110011001100110011001101001011010011001011010010110,
64'b1111111111111111000000000000000010100101101001010101101001011010,
64'b0011001111001100001100111100110011111111111111110000000000000000,
64'b0000000011111111111111110000000001101001011010011001011010010110,
64'b0000000000000000000000000000000000001111111100000000111111110000,
64'b0101101001011010010110100101101001010101010101011010101010101010,
64'b0011110011000011110000110011110011110000111100001111000011110000,
64'b0000000011111111111111110000000010100101101001010101101001011010,
64'b0110011001100110011001100110011011000011110000110011110000111100,
64'b0011001111001100001100111100110000110011001100111100110011001100,
64'b1111000000001111000011111111000010011001011001101001100101100110,
64'b1100110000110011001100111100110011000011001111001100001100111100,
64'b1100110011001100110011001100110010011001011001101001100101100110,
64'b0101101001011010010110100101101011110000000011110000111111110000,
64'b0101101001011010010110100101101010100101010110101010010101011010,
64'b1001100101100110100110010110011001011010010110100101101001011010,
64'b1010101001010101010101011010101010101010010101010101010110101010,
64'b1001011010010110100101101001011011111111000000001111111100000000,
64'b1100001100111100110000110011110001100110011001100110011001100110,
64'b1100110011001100110011001100110001010101101010100101010110101010,
64'b0101010110101010010101011010101000110011110011000011001111001100,
64'b1111000011110000111100001111000010100101010110101010010101011010,
64'b0011110011000011110000110011110001011010010110100101101001011010,
64'b1111000011110000111100001111000001101001011010011001011010010110,
64'b0110100110010110011010011001011011110000000011110000111111110000,
64'b1001011010010110100101101001011011000011110000110011110000111100,
64'b0110100110010110011010011001011000000000111111111111111100000000,
64'b0110100110010110011010011001011001100110100110011001100101100110,
64'b0101101010100101101001010101101000110011110011000011001111001100,
64'b1001100101100110100110010110011000110011001100111100110011001100,
64'b1111111100000000111111110000000010101010101010101010101010101010,
64'b0000000011111111111111110000000000111100001111000011110000111100,
64'b1100110000110011001100111100110000110011001100111100110011001100,
64'b0011001111001100001100111100110000001111000011111111000011110000,
64'b1001100101100110100110010110011011001100001100110011001111001100,
64'b1100001111000011001111000011110000110011110011000011001111001100,
64'b1010010110100101010110100101101011000011001111001100001100111100,
64'b1111000011110000111100001111000010101010010101010101010110101010,
64'b0000111111110000000011111111000010100101010110101010010101011010,
64'b0110011010011001100110010110011001010101010101011010101010101010,
64'b0110011010011001100110010110011001101001011010011001011010010110,
64'b0101010101010101101010101010101010100101101001010101101001011010,
64'b1100001100111100110000110011110011110000111100001111000011110000,
64'b1001011010010110100101101001011001100110011001100110011001100110,
64'b0101010101010101101010101010101000001111111100000000111111110000,
64'b1010010110100101010110100101101011110000111100001111000011110000,
64'b1010010110100101010110100101101001010101101010100101010110101010,
64'b1100001111000011001111000011110010100101101001010101101001011010,
64'b0000111111110000000011111111000010100101101001010101101001011010,
64'b1001100101100110100110010110011011110000000011110000111111110000,
64'b0101010110101010010101011010101000110011001100111100110011001100,
64'b0000000011111111111111110000000001100110100110011001100101100110,
64'b1100001111000011001111000011110011001100110011001100110011001100,
64'b0110100101101001100101101001011001101001100101100110100110010110,
64'b0110011001100110011001100110011010011001011001101001100101100110,
64'b0101101010100101101001010101101001010101101010100101010110101010,
64'b1100001100111100110000110011110000111100001111000011110000111100,
64'b0011110000111100001111000011110000000000111111111111111100000000,
64'b1010010110100101010110100101101011111111000000001111111100000000,
64'b1001100110011001011001100110011000110011001100111100110011001100,
64'b1100001100111100110000110011110000110011110011000011001111001100,
64'b1001100110011001011001100110011010011001011001101001100101100110,
64'b0011001111001100001100111100110010101010010101010101010110101010,
64'b1111111100000000111111110000000001011010010110100101101001011010,
64'b0011001100110011110011001100110001101001011010011001011010010110,
64'b1111111100000000111111110000000001011010010110100101101001011010,
64'b0011001111001100001100111100110000111100110000111100001100111100,
64'b0000111111110000000011111111000011000011110000110011110000111100,
64'b0110011001100110011001100110011000110011001100111100110011001100,
64'b0011001111001100001100111100110000001111111100000000111111110000,
64'b0101010110101010010101011010101001010101010101011010101010101010,
64'b0000111100001111111100001111000001010101010101011010101010101010,
64'b1001011001101001011010011001011011110000111100001111000011110000,
64'b0011110011000011110000110011110010100101101001010101101001011010,
64'b0000111111110000000011111111000011000011110000110011110000111100,
64'b0101010110101010010101011010101000110011001100111100110011001100,
64'b0011001111001100001100111100110010011001011001101001100101100110,
64'b0011110000111100001111000011110011000011001111001100001100111100,
64'b0000111100001111111100001111000010011001011001101001100101100110,
64'b0101010101010101101010101010101011110000000011110000111111110000,
64'b1001100110011001011001100110011010100101010110101010010101011010,
64'b1001011001101001011010011001011001011010010110100101101001011010,
64'b0110011001100110011001100110011001010101101010100101010110101010,
64'b1001100110011001011001100110011000111100001111000011110000111100,
64'b1111111100000000111111110000000001011010101001011010010101011010,
64'b1001011001101001011010011001011001010101010101011010101010101010,
64'b0101101010100101101001010101101001010101101010100101010110101010,
64'b1010101001010101010101011010101010010110100101101001011010010110,
64'b0011001100110011110011001100110010101010010101010101010110101010,
64'b0000111100001111111100001111000010100101010110101010010101011010,
64'b0000111111110000000011111111000000111100110000111100001100111100,
64'b1111111100000000111111110000000010011001100110010110011001100110,
64'b0110011001100110011001100110011001011010101001011010010101011010,
64'b1001011010010110100101101001011011111111111111110000000000000000,
64'b1001011001101001011010011001011010011001100110010110011001100110,
64'b1001011010010110100101101001011001011010010110100101101001011010,
64'b0110011001100110011001100110011001010101101010100101010110101010,
64'b0110100110010110011010011001011011110000111100001111000011110000,
64'b0011110000111100001111000011110001100110100110011001100101100110,
64'b0000000011111111111111110000000011111111111111110000000000000000,
64'b1010101001010101010101011010101011110000111100001111000011110000,
64'b1010101001010101010101011010101011000011001111001100001100111100,
64'b1001100110011001011001100110011010101010101010101010101010101010,
64'b0110011010011001100110010110011000111100110000111100001100111100,
64'b1010010110100101010110100101101011001100110011001100110011001100,
64'b0110011001100110011001100110011000111100110000111100001100111100,
64'b0101101001011010010110100101101000110011110011000011001111001100,
64'b1001011010010110100101101001011000111100110000111100001100111100,
64'b1111111100000000111111110000000000001111111100000000111111110000,
64'b1100110011001100110011001100110000110011001100111100110011001100,
64'b0000000000000000000000000000000011111111000000001111111100000000,
64'b0000111100001111111100001111000011000011110000110011110000111100,
64'b1001100110011001011001100110011010101010101010101010101010101010,
64'b1010101001010101010101011010101001010101101010100101010110101010,
64'b0110100110010110011010011001011011110000000011110000111111110000,
64'b0101101010100101101001010101101011001100110011001100110011001100,
64'b1010010110100101010110100101101011110000000011110000111111110000,
64'b1100001100111100110000110011110001011010010110100101101001011010,
64'b1100110011001100110011001100110011110000000011110000111111110000,
64'b1010101010101010101010101010101010100101101001010101101001011010,
64'b0110100101101001100101101001011011110000000011110000111111110000,
64'b1001011010010110100101101001011001010101101010100101010110101010,
64'b0101101001011010010110100101101001011010010110100101101001011010,
64'b0000000000000000000000000000000001010101010101011010101010101010,
64'b1111111100000000111111110000000000001111111100000000111111110000,
64'b1001011010010110100101101001011001100110011001100110011001100110,
64'b1001100110011001011001100110011000110011001100111100110011001100,
64'b1001011001101001011010011001011000000000111111111111111100000000,
64'b1100110000110011001100111100110001011010010110100101101001011010,
64'b1001100101100110100110010110011000000000111111111111111100000000,
64'b0101101010100101101001010101101010011001011001101001100101100110,
64'b1111000011110000111100001111000000000000111111111111111100000000,
64'b1100110011001100110011001100110010011001011001101001100101100110,
64'b1100001100111100110000110011110010101010010101010101010110101010,
64'b0110100110010110011010011001011001100110011001100110011001100110,
64'b1100001100111100110000110011110001101001100101100110100110010110,
64'b0011110011000011110000110011110011110000000011110000111111110000,
64'b1111111100000000111111110000000010101010101010101010101010101010,
64'b1010010101011010101001010101101001011010010110100101101001011010,
64'b0000111111110000000011111111000011000011001111001100001100111100,
64'b0110011001100110011001100110011010100101010110101010010101011010,
64'b0110100110010110011010011001011001010101010101011010101010101010,
64'b1010010110100101010110100101101000110011001100111100110011001100,
64'b1001011001101001011010011001011000110011001100111100110011001100,
64'b0000111111110000000011111111000010100101101001010101101001011010,
64'b0110100110010110011010011001011011110000000011110000111111110000,
64'b0101101001011010010110100101101010011001011001101001100101100110,
64'b0101010110101010010101011010101000000000000000000000000000000000,
64'b0000000011111111111111110000000000111100110000111100001100111100,
64'b1100110011001100110011001100110000000000111111111111111100000000,
64'b0101010110101010010101011010101001100110011001100110011001100110,
64'b1010101001010101010101011010101000110011110011000011001111001100,
64'b0011001100110011110011001100110011110000000011110000111111110000,
64'b1100110000110011001100111100110011001100001100110011001111001100,
64'b1111000011110000111100001111000011001100110011001100110011001100,
64'b1111111100000000111111110000000001011010010110100101101001011010,
64'b1100110000110011001100111100110001011010010110100101101001011010,
64'b1111000000001111000011111111000010011001011001101001100101100110,
64'b1010010110100101010110100101101010101010010101010101010110101010,
64'b1001100110011001011001100110011001101001011010011001011010010110,
64'b0101101001011010010110100101101000000000000000000000000000000000,
64'b1010010110100101010110100101101011110000000011110000111111110000,
64'b0110011010011001100110010110011001010101010101011010101010101010,
64'b0011001111001100001100111100110010010110100101101001011010010110,
64'b0101010101010101101010101010101000001111000011111111000011110000,
64'b0110100110010110011010011001011000000000111111111111111100000000,
64'b0101010110101010010101011010101010100101101001010101101001011010,
64'b1001100110011001011001100110011001011010010110100101101001011010,
64'b0011001100110011110011001100110000110011110011000011001111001100,
64'b0101010101010101101010101010101000110011110011000011001111001100,
64'b1111000000001111000011111111000011000011110000110011110000111100,
64'b0000000000000000000000000000000000110011001100111100110011001100,
64'b0011110011000011110000110011110001101001100101100110100110010110,
64'b0000111111110000000011111111000010101010101010101010101010101010,
64'b0011001111001100001100111100110000000000111111111111111100000000,
64'b0110100101101001100101101001011001100110011001100110011001100110,
64'b1010010110100101010110100101101001101001100101100110100110010110,
64'b1100110011001100110011001100110011111111000000001111111100000000,
64'b1001011001101001011010011001011001010101010101011010101010101010,
64'b0011001100110011110011001100110010011001011001101001100101100110,
64'b0011110000111100001111000011110010011001011001101001100101100110,
64'b0101101001011010010110100101101000001111000011111111000011110000,
64'b0110011001100110011001100110011000001111000011111111000011110000,
64'b1010101001010101010101011010101000001111111100000000111111110000,
64'b1010101010101010101010101010101001011010010110100101101001011010,
64'b1111000000001111000011111111000010010110011010010110100110010110,
64'b0101010110101010010101011010101011001100110011001100110011001100,
64'b1010010110100101010110100101101001010101010101011010101010101010,
64'b1100001100111100110000110011110010010110100101101001011010010110,
64'b1001100101100110100110010110011000111100110000111100001100111100,
64'b0101101001011010010110100101101011111111111111110000000000000000,
64'b0011110011000011110000110011110011001100110011001100110011001100,
64'b0101101001011010010110100101101001101001011010011001011010010110,
64'b1010010101011010101001010101101011000011110000110011110000111100,
64'b0011001111001100001100111100110011111111000000001111111100000000,
64'b0011110000111100001111000011110001010101101010100101010110101010,
64'b0011001100110011110011001100110010101010010101010101010110101010,
64'b0110011001100110011001100110011000110011110011000011001111001100,
64'b0000000011111111111111110000000000111100110000111100001100111100,
64'b0110011001100110011001100110011001011010010110100101101001011010,
64'b0011001111001100001100111100110011001100110011001100110011001100,
64'b0101101010100101101001010101101001101001100101100110100110010110,
64'b1100001111000011001111000011110011110000000011110000111111110000,
64'b0011001111001100001100111100110010101010101010101010101010101010,
64'b1111000000001111000011111111000001011010010110100101101001011010,
64'b1001100101100110100110010110011011000011001111001100001100111100,
64'b1100110000110011001100111100110010100101010110101010010101011010,
64'b0000111100001111111100001111000001010101010101011010101010101010,
64'b0000111111110000000011111111000000110011001100111100110011001100,
64'b1111000011110000111100001111000000110011001100111100110011001100,
64'b1001011010010110100101101001011010100101101001010101101001011010,
64'b1111111111111111000000000000000011110000000011110000111111110000,
64'b1001011010010110100101101001011010011001011001101001100101100110,
64'b1010101010101010101010101010101001011010101001011010010101011010,
64'b0011110011000011110000110011110011000011001111001100001100111100,
64'b0011110011000011110000110011110001100110011001100110011001100110,
64'b0110100101101001100101101001011000001111000011111111000011110000,
64'b1001100110011001011001100110011001100110100110011001100101100110,
64'b1010010101011010101001010101101000110011110011000011001111001100,
64'b1010101001010101010101011010101000111100001111000011110000111100,
64'b0011110011000011110000110011110011110000111100001111000011110000,
64'b0101101010100101101001010101101000001111111100000000111111110000,
64'b1100001111000011001111000011110001101001100101100110100110010110,
64'b1100001111000011001111000011110001101001100101100110100110010110,
64'b1111111100000000111111110000000000000000111111111111111100000000,
64'b1100110011001100110011001100110000111100001111000011110000111100,
64'b0110011001100110011001100110011001100110100110011001100101100110,
64'b1100110011001100110011001100110001011010101001011010010101011010,
64'b0110011001100110011001100110011000111100001111000011110000111100,
64'b0000000011111111111111110000000011111111000000001111111100000000,
64'b0000111100001111111100001111000001101001011010011001011010010110,
64'b1100001111000011001111000011110010100101101001010101101001011010,
64'b1001100101100110100110010110011000001111111100000000111111110000,
64'b0110011001100110011001100110011011111111000000001111111100000000,
64'b0011110000111100001111000011110000000000111111111111111100000000,
64'b0110011010011001100110010110011000111100110000111100001100111100,
64'b0110011010011001100110010110011000111100110000111100001100111100,
64'b1010101001010101010101011010101011111111111111110000000000000000,
64'b0011110000111100001111000011110010100101010110101010010101011010,
64'b0011110000111100001111000011110011000011110000110011110000111100,
64'b1100110000110011001100111100110001100110100110011001100101100110,
64'b0000000011111111111111110000000010100101010110101010010101011010,
64'b1001011010010110100101101001011011111111111111110000000000000000,
64'b1100110000110011001100111100110011000011001111001100001100111100,
64'b0000000000000000000000000000000010011001011001101001100101100110,
64'b1100001100111100110000110011110010101010010101010101010110101010,
64'b0000000011111111111111110000000011111111111111110000000000000000,
64'b0101010101010101101010101010101011111111111111110000000000000000,
64'b0000000000000000000000000000000001011010101001011010010101011010,
64'b1010101010101010101010101010101001011010101001011010010101011010,
64'b0110011010011001100110010110011010101010101010101010101010101010,
64'b0110100110010110011010011001011010011001011001101001100101100110,
64'b0000111111110000000011111111000000001111111100000000111111110000,
64'b0000111100001111111100001111000001101001011010011001011010010110,
64'b0101010101010101101010101010101001100110100110011001100101100110,
64'b0110100110010110011010011001011000000000000000000000000000000000,
64'b0000111100001111111100001111000001011010101001011010010101011010,
64'b1010101010101010101010101010101011000011110000110011110000111100,
64'b1111000000001111000011111111000000110011001100111100110011001100,
64'b1111111111111111000000000000000010101010101010101010101010101010,
64'b0110011001100110011001100110011010101010101010101010101010101010,
64'b1010101010101010101010101010101001100110100110011001100101100110,
64'b1100110011001100110011001100110001100110100110011001100101100110,
64'b1100001111000011001111000011110001100110011001100110011001100110,
64'b0110100110010110011010011001011000111100001111000011110000111100,
64'b0000000011111111111111110000000000000000111111111111111100000000,
64'b1100001111000011001111000011110011000011001111001100001100111100,
64'b0101101010100101101001010101101001101001011010011001011010010110,
64'b1111111100000000111111110000000010101010101010101010101010101010,
64'b0110011010011001100110010110011011001100001100110011001111001100,
64'b1100001100111100110000110011110010100101010110101010010101011010,
64'b1010101010101010101010101010101001011010010110100101101001011010,
64'b1001011001101001011010011001011001100110011001100110011001100110,
64'b1100110000110011001100111100110011001100110011001100110011001100,
64'b0000111100001111111100001111000011000011110000110011110000111100,
64'b0011001100110011110011001100110001101001011010011001011010010110,
64'b1111000011110000111100001111000010010110100101101001011010010110,
64'b1010010101011010101001010101101000001111111100000000111111110000,
64'b1111111111111111000000000000000001010101010101011010101010101010,
64'b1001100110011001011001100110011001011010101001011010010101011010,
64'b0101101001011010010110100101101011000011001111001100001100111100,
64'b0011110000111100001111000011110001100110011001100110011001100110,
64'b0101101001011010010110100101101000001111000011111111000011110000,
64'b1111111111111111000000000000000001100110100110011001100101100110,
64'b0110011010011001100110010110011000110011110011000011001111001100,
64'b0000000000000000000000000000000000111100001111000011110000111100,
64'b1111111100000000111111110000000011110000111100001111000011110000,
64'b1001011001101001011010011001011000001111111100000000111111110000,
64'b1001100110011001011001100110011001101001100101100110100110010110,
64'b1010101010101010101010101010101001101001100101100110100110010110,
64'b1111111100000000111111110000000011111111000000001111111100000000,
64'b0000000000000000000000000000000011001100110011001100110011001100,
64'b1001011010010110100101101001011001011010010110100101101001011010,
64'b1001100101100110100110010110011001100110011001100110011001100110,
64'b0000111111110000000011111111000001010101010101011010101010101010,
64'b0011001111001100001100111100110001100110100110011001100101100110,
64'b0000000000000000000000000000000011001100001100110011001111001100,
64'b0110100101101001100101101001011000001111111100000000111111110000,
64'b1010101010101010101010101010101000110011001100111100110011001100,
64'b1111111111111111000000000000000010100101101001010101101001011010,
64'b0011110011000011110000110011110011000011001111001100001100111100,
64'b1001011010010110100101101001011011111111000000001111111100000000,
64'b0110011001100110011001100110011011000011110000110011110000111100,
64'b0000000000000000000000000000000011001100110011001100110011001100,
64'b1010101010101010101010101010101001011010010110100101101001011010,
64'b1111111111111111000000000000000000001111000011111111000011110000,
64'b1111111100000000111111110000000000000000111111111111111100000000,
64'b0110100110010110011010011001011010100101101001010101101001011010,
64'b1001011010010110100101101001011011110000111100001111000011110000,
64'b1010010101011010101001010101101000000000111111111111111100000000,
64'b0110100101101001100101101001011000000000000000000000000000000000,
64'b0101101010100101101001010101101011001100001100110011001111001100,
64'b0101101010100101101001010101101011000011110000110011110000111100,
64'b1001100101100110100110010110011010011001011001101001100101100110,
64'b1010101001010101010101011010101000111100001111000011110000111100,
64'b1100001100111100110000110011110011110000111100001111000011110000,
64'b1100110011001100110011001100110010010110100101101001011010010110,
64'b1100110011001100110011001100110010011001011001101001100101100110,
64'b0011110011000011110000110011110011111111000000001111111100000000,
64'b0110100110010110011010011001011001010101010101011010101010101010,
64'b0101010110101010010101011010101010011001011001101001100101100110,
64'b0101101010100101101001010101101001010101101010100101010110101010,
64'b0110100101101001100101101001011011111111111111110000000000000000,
64'b0110100101101001100101101001011010101010101010101010101010101010,
64'b0101101001011010010110100101101000001111000011111111000011110000,
64'b0011110000111100001111000011110010100101010110101010010101011010,
64'b1010101010101010101010101010101001101001011010011001011010010110,
64'b1111000011110000111100001111000000001111111100000000111111110000,
64'b1010010110100101010110100101101011111111000000001111111100000000,
64'b0011110000111100001111000011110011000011001111001100001100111100,
64'b1111000011110000111100001111000001101001011010011001011010010110,
64'b1111000000001111000011111111000011111111111111110000000000000000,
64'b1001011001101001011010011001011011001100110011001100110011001100,
64'b0011001100110011110011001100110001101001011010011001011010010110,
64'b1100110000110011001100111100110000110011001100111100110011001100,
64'b0110100110010110011010011001011000000000000000000000000000000000,
64'b0110100110010110011010011001011001100110011001100110011001100110,
64'b1001100101100110100110010110011011111111000000001111111100000000,
64'b0000111111110000000011111111000001100110100110011001100101100110,
64'b1100110011001100110011001100110011000011001111001100001100111100,
64'b1111111100000000111111110000000010101010010101010101010110101010,
64'b0011001111001100001100111100110011111111111111110000000000000000,
64'b1010010101011010101001010101101000001111111100000000111111110000,
64'b1111111100000000111111110000000001101001100101100110100110010110,
64'b0011110000111100001111000011110010010110011010010110100110010110,
64'b1010101010101010101010101010101001100110100110011001100101100110,
64'b0011001100110011110011001100110010101010010101010101010110101010,
64'b0011110000111100001111000011110011000011110000110011110000111100,
64'b0011001100110011110011001100110000001111111100000000111111110000,
64'b1001011010010110100101101001011010010110011010010110100110010110,
64'b1111111100000000111111110000000011000011001111001100001100111100,
64'b0101101001011010010110100101101010011001011001101001100101100110,
64'b0011001100110011110011001100110010011001011001101001100101100110,
64'b0011110000111100001111000011110011110000111100001111000011110000,
64'b1111000000001111000011111111000001010101101010100101010110101010,
64'b1111111100000000111111110000000010011001011001101001100101100110,
64'b1111111111111111000000000000000000111100110000111100001100111100,
64'b0011001100110011110011001100110000111100110000111100001100111100,
64'b1111000000001111000011111111000001101001011010011001011010010110,
64'b1001100110011001011001100110011010011001100110010110011001100110,
64'b0011110011000011110000110011110010100101010110101010010101011010,
64'b0101010110101010010101011010101010101010010101010101010110101010,
64'b1100001111000011001111000011110000111100110000111100001100111100,
64'b1100001100111100110000110011110001011010101001011010010101011010,
64'b0110100101101001100101101001011011000011110000110011110000111100,
64'b0011001100110011110011001100110011000011110000110011110000111100,
64'b0110011010011001100110010110011011111111000000001111111100000000,
64'b1111111111111111000000000000000000110011001100111100110011001100,
64'b0110011001100110011001100110011000111100001111000011110000111100,
64'b1010101010101010101010101010101011110000000011110000111111110000,
64'b0110011010011001100110010110011001011010101001011010010101011010,
64'b1001011010010110100101101001011001101001100101100110100110010110,
64'b1111111111111111000000000000000010010110100101101001011010010110,
64'b1100001100111100110000110011110001100110100110011001100101100110,
64'b0011110011000011110000110011110000110011001100111100110011001100,
64'b1010010110100101010110100101101001011010101001011010010101011010,
64'b0110011001100110011001100110011001100110100110011001100101100110,
64'b1001100110011001011001100110011010100101010110101010010101011010,
64'b1001100110011001011001100110011010100101010110101010010101011010,
64'b1010101010101010101010101010101001010101010101011010101010101010,
64'b0101010110101010010101011010101011110000111100001111000011110000,
64'b0101101001011010010110100101101010100101010110101010010101011010,
64'b0110011001100110011001100110011000000000111111111111111100000000,
64'b1100001111000011001111000011110001100110100110011001100101100110,
64'b0110100110010110011010011001011010010110011010010110100110010110,
64'b0000000000000000000000000000000011000011001111001100001100111100,
64'b0101101010100101101001010101101011000011110000110011110000111100,
64'b1111000000001111000011111111000001011010010110100101101001011010,
64'b1001100101100110100110010110011001100110100110011001100101100110,
64'b1001011010010110100101101001011001101001011010011001011010010110,
64'b0011110000111100001111000011110001100110100110011001100101100110,
64'b1001011010010110100101101001011011001100001100110011001111001100,
64'b0110011001100110011001100110011011001100110011001100110011001100,
64'b0011001100110011110011001100110001010101101010100101010110101010,
64'b0011001111001100001100111100110000110011110011000011001111001100,
64'b1001011010010110100101101001011011111111111111110000000000000000,
64'b0000111111110000000011111111000001101001011010011001011010010110,
64'b1001011001101001011010011001011010010110011010010110100110010110,
64'b0000000000000000000000000000000001011010101001011010010101011010,
64'b1100110000110011001100111100110000001111111100000000111111110000,
64'b1010101001010101010101011010101010011001011001101001100101100110,
64'b0110100101101001100101101001011011000011110000110011110000111100,
64'b1100001100111100110000110011110001101001100101100110100110010110,
64'b0000111111110000000011111111000001101001011010011001011010010110,
64'b1100001100111100110000110011110010100101101001010101101001011010,
64'b0011110000111100001111000011110001011010010110100101101001011010,
64'b1111000011110000111100001111000000110011001100111100110011001100,
64'b0101101001011010010110100101101011110000111100001111000011110000,
64'b1100001100111100110000110011110000000000000000000000000000000000,
64'b0000000011111111111111110000000001101001100101100110100110010110,
64'b0011110011000011110000110011110010010110011010010110100110010110,
64'b1010101010101010101010101010101001100110100110011001100101100110,
64'b0000111100001111111100001111000010101010010101010101010110101010,
64'b1001100110011001011001100110011011000011110000110011110000111100,
64'b0110100110010110011010011001011000001111111100000000111111110000,
64'b0101101010100101101001010101101010010110011010010110100110010110,
64'b0000000011111111111111110000000011000011001111001100001100111100,
64'b1111000000001111000011111111000010011001011001101001100101100110,
64'b0000111111110000000011111111000010011001011001101001100101100110,
64'b1111111100000000111111110000000011110000111100001111000011110000,
64'b0011001111001100001100111100110001010101101010100101010110101010,
64'b1010010101011010101001010101101000000000111111111111111100000000,
64'b1010010101011010101001010101101001101001011010011001011010010110,
64'b1100110000110011001100111100110010010110100101101001011010010110,
64'b0110100110010110011010011001011010010110100101101001011010010110,
64'b0110100101101001100101101001011010010110011010010110100110010110,
64'b1010101001010101010101011010101011110000111100001111000011110000,
64'b0101010101010101101010101010101001011010010110100101101001011010,
64'b0000000011111111111111110000000010010110100101101001011010010110,
64'b1010101010101010101010101010101000110011110011000011001111001100,
64'b1010010101011010101001010101101011110000111100001111000011110000,
64'b0101101001011010010110100101101010100101010110101010010101011010,
64'b0101101001011010010110100101101010101010010101010101010110101010,
64'b0101101001011010010110100101101010100101010110101010010101011010,
64'b0110100101101001100101101001011011111111111111110000000000000000,
64'b0110100101101001100101101001011001101001100101100110100110010110,
64'b1100001100111100110000110011110001101001100101100110100110010110,
64'b1111111111111111000000000000000011000011001111001100001100111100,
64'b1010101001010101010101011010101000111100110000111100001100111100,
64'b0011001111001100001100111100110001010101101010100101010110101010,
64'b0011001100110011110011001100110000110011110011000011001111001100,
64'b0101010110101010010101011010101011000011001111001100001100111100,
64'b1100110011001100110011001100110000001111000011111111000011110000,
64'b0110100101101001100101101001011011111111000000001111111100000000,
64'b0110100110010110011010011001011011001100001100110011001111001100,
64'b0110100110010110011010011001011000110011001100111100110011001100,
64'b0110100110010110011010011001011010011001011001101001100101100110,
64'b0110011001100110011001100110011010101010101010101010101010101010,
64'b1100110011001100110011001100110010010110011010010110100110010110,
64'b1001011010010110100101101001011000111100110000111100001100111100,
64'b0110100110010110011010011001011011110000000011110000111111110000,
64'b1111000011110000111100001111000011110000000011110000111111110000,
64'b0000111111110000000011111111000010011001100110010110011001100110,
64'b1010010110100101010110100101101000001111000011111111000011110000,
64'b1001100101100110100110010110011011110000000011110000111111110000,
64'b0101101001011010010110100101101011111111000000001111111100000000,
64'b0110011001100110011001100110011001010101010101011010101010101010,
64'b1100110000110011001100111100110000001111000011111111000011110000,
64'b0110011010011001100110010110011001011010010110100101101001011010,
64'b1001100101100110100110010110011010010110100101101001011010010110,
64'b1001011010010110100101101001011001100110011001100110011001100110,
64'b1111000011110000111100001111000000111100110000111100001100111100,
64'b1100001100111100110000110011110001011010101001011010010101011010,
64'b0011110011000011110000110011110010101010010101010101010110101010,
64'b1111111100000000111111110000000010101010010101010101010110101010,
64'b0000000011111111111111110000000010010110100101101001011010010110,
64'b0011001111001100001100111100110001010101101010100101010110101010,
64'b0110100101101001100101101001011010101010010101010101010110101010,
64'b0011001111001100001100111100110001010101010101011010101010101010,
64'b0011110000111100001111000011110011001100110011001100110011001100,
64'b0000111100001111111100001111000001010101101010100101010110101010,
64'b0110100101101001100101101001011010011001011001101001100101100110,
64'b1001011010010110100101101001011011000011001111001100001100111100,
64'b1100110011001100110011001100110000111100001111000011110000111100,
64'b0101101001011010010110100101101011110000000011110000111111110000,
64'b0011110000111100001111000011110001100110100110011001100101100110,
64'b1001100110011001011001100110011010011001100110010110011001100110,
64'b0011110000111100001111000011110010011001100110010110011001100110,
64'b0101010110101010010101011010101001101001100101100110100110010110,
64'b1111000011110000111100001111000000110011001100111100110011001100,
64'b1100001111000011001111000011110000110011001100111100110011001100,
64'b0000111100001111111100001111000001100110011001100110011001100110,
64'b1010101010101010101010101010101001011010010110100101101001011010,
64'b1010010101011010101001010101101000110011001100111100110011001100,
64'b0011001111001100001100111100110011000011110000110011110000111100,
64'b0011001111001100001100111100110000001111111100000000111111110000,
64'b1111111100000000111111110000000010100101010110101010010101011010,
64'b1001011010010110100101101001011000000000111111111111111100000000,
64'b1100001111000011001111000011110001101001011010011001011010010110,
64'b0101010110101010010101011010101010010110100101101001011010010110,
64'b1100110000110011001100111100110010010110100101101001011010010110,
64'b1001100101100110100110010110011010010110011010010110100110010110,
64'b1010101001010101010101011010101011110000111100001111000011110000,
64'b0000111100001111111100001111000001011010010110100101101001011010,
64'b1111111100000000111111110000000010010110100101101001011010010110,
64'b1100001100111100110000110011110000110011110011000011001111001100,
64'b1001011001101001011010011001011011110000111100001111000011110000,
64'b0101010101010101101010101010101010100101010110101010010101011010,
64'b1010101010101010101010101010101001010101101010100101010110101010,
64'b0101010101010101101010101010101011000011110000110011110000111100,
64'b1100001100111100110000110011110001011010101001011010010101011010,
64'b0000111111110000000011111111000010100101101001010101101001011010,
64'b1001100110011001011001100110011000000000000000000000000000000000,
64'b0000111100001111111100001111000010101010010101010101010110101010,
64'b0110100101101001100101101001011010010110100101101001011010010110,
64'b0011001100110011110011001100110000000000111111111111111100000000,
64'b0101010110101010010101011010101000110011001100111100110011001100,
64'b0101010101010101101010101010101001101001100101100110100110010110,
64'b1111000000001111000011111111000010101010010101010101010110101010,
64'b0011110011000011110000110011110010100101010110101010010101011010,
64'b0110011001100110011001100110011010010110011010010110100110010110,
64'b0110011001100110011001100110011010010110100101101001011010010110,
64'b0110100110010110011010011001011010101010101010101010101010101010,
64'b1111111111111111000000000000000011000011110000110011110000111100,
64'b1100110011001100110011001100110001010101010101011010101010101010,
64'b0101010110101010010101011010101011000011001111001100001100111100,
64'b0011110011000011110000110011110001011010010110100101101001011010,
64'b1100001111000011001111000011110011000011110000110011110000111100,
64'b0000111100001111111100001111000010101010101010101010101010101010,
64'b1001100101100110100110010110011001011010101001011010010101011010,
64'b0110011001100110011001100110011000111100110000111100001100111100,
64'b0000111100001111111100001111000010010110011010010110100110010110,
64'b0000000011111111111111110000000000111100110000111100001100111100,
64'b1100110011001100110011001100110001100110100110011001100101100110,
64'b0110011001100110011001100110011000110011110011000011001111001100,
64'b1001100110011001011001100110011011001100110011001100110011001100,
64'b1010010101011010101001010101101000001111111100000000111111110000,
64'b1001011001101001011010011001011001100110011001100110011001100110,
64'b0101101010100101101001010101101001011010101001011010010101011010,
64'b1001100101100110100110010110011000110011110011000011001111001100,
64'b0000111100001111111100001111000000001111111100000000111111110000,
64'b0000000011111111111111110000000001100110011001100110011001100110,
64'b0110100110010110011010011001011011001100001100110011001111001100,
64'b1001011010010110100101101001011001011010101001011010010101011010,
64'b0101101001011010010110100101101010010110011010010110100110010110,
64'b0000111100001111111100001111000001011010101001011010010101011010,
64'b0000000000000000000000000000000001101001011010011001011010010110,
64'b0110011001100110011001100110011001011010010110100101101001011010,
64'b0011110000111100001111000011110001011010010110100101101001011010,
64'b0110011010011001100110010110011000000000111111111111111100000000,
64'b0011110011000011110000110011110000111100001111000011110000111100,
64'b0110011010011001100110010110011011001100001100110011001111001100,
64'b0110100101101001100101101001011010100101101001010101101001011010,
64'b1111111100000000111111110000000000000000111111111111111100000000,
64'b0101010101010101101010101010101000111100001111000011110000111100,
64'b1001011001101001011010011001011000001111000011111111000011110000,
64'b1100001100111100110000110011110001100110100110011001100101100110,
64'b0011001111001100001100111100110010010110011010010110100110010110,
64'b1111111100000000111111110000000001100110100110011001100101100110,
64'b1010101010101010101010101010101001101001100101100110100110010110,
64'b0011110000111100001111000011110010011001011001101001100101100110,
64'b0000000000000000000000000000000000111100001111000011110000111100,
64'b0110011010011001100110010110011001011010101001011010010101011010,
64'b1001011010010110100101101001011001101001011010011001011010010110,
64'b0000000011111111111111110000000001100110100110011001100101100110,
64'b0000000011111111111111110000000011110000000011110000111111110000,
64'b1111111100000000111111110000000011111111000000001111111100000000,
64'b1001100110011001011001100110011011110000000011110000111111110000,
64'b1001011010010110100101101001011011111111111111110000000000000000,
64'b1111000000001111000011111111000011000011110000110011110000111100,
64'b1010101001010101010101011010101000110011001100111100110011001100,
64'b1010010110100101010110100101101000110011001100111100110011001100,
64'b1001011010010110100101101001011011001100001100110011001111001100,
64'b0101010110101010010101011010101001100110011001100110011001100110,
64'b0000111111110000000011111111000010100101010110101010010101011010,
64'b0110011010011001100110010110011011001100001100110011001111001100,
64'b1010010110100101010110100101101001101001100101100110100110010110,
64'b1001011001101001011010011001011001101001011010011001011010010110,
64'b0011110000111100001111000011110010101010010101010101010110101010,
64'b1111111100000000111111110000000001010101010101011010101010101010,
64'b0110100101101001100101101001011000000000111111111111111100000000,
64'b0110100101101001100101101001011010101010101010101010101010101010,
64'b1010101001010101010101011010101010100101010110101010010101011010,
64'b0011110011000011110000110011110001011010010110100101101001011010,
64'b1100001100111100110000110011110001011010010110100101101001011010,
64'b0011001111001100001100111100110010100101101001010101101001011010,
64'b1001011010010110100101101001011010010110100101101001011010010110,
64'b1010010110100101010110100101101011001100001100110011001111001100,
64'b0110011010011001100110010110011000001111000011111111000011110000,
64'b0101010101010101101010101010101010010110011010010110100110010110,
64'b1111111111111111000000000000000011000011001111001100001100111100,
64'b1100110000110011001100111100110010011001100110010110011001100110,
64'b0101010110101010010101011010101001100110011001100110011001100110,
64'b1001011001101001011010011001011001010101010101011010101010101010,
64'b0110100101101001100101101001011001100110011001100110011001100110,
64'b0011001100110011110011001100110011001100001100110011001111001100,
64'b1111111111111111000000000000000000110011110011000011001111001100,
64'b0000000011111111111111110000000000110011110011000011001111001100,
64'b0101010101010101101010101010101000110011110011000011001111001100,
64'b1001100101100110100110010110011001101001100101100110100110010110,
64'b0011001111001100001100111100110010100101101001010101101001011010,
64'b0110100101101001100101101001011001010101101010100101010110101010,
64'b0110011001100110011001100110011010010110011010010110100110010110,
64'b1010101010101010101010101010101001011010101001011010010101011010,
64'b1010010110100101010110100101101000111100001111000011110000111100,
64'b1001100110011001011001100110011010010110100101101001011010010110,
64'b0011110011000011110000110011110011001100110011001100110011001100,
64'b0110100110010110011010011001011010010110100101101001011010010110,
64'b0101101001011010010110100101101000001111000011111111000011110000,
64'b1010101010101010101010101010101010100101101001010101101001011010,
64'b0101010101010101101010101010101000001111000011111111000011110000,
64'b0110011001100110011001100110011000001111000011111111000011110000,
64'b1001011010010110100101101001011011000011001111001100001100111100,
64'b1010010110100101010110100101101010011001011001101001100101100110,
64'b1100001100111100110000110011110010011001100110010110011001100110,
64'b1001011010010110100101101001011000111100110000111100001100111100,
64'b1100110011001100110011001100110001100110100110011001100101100110,
64'b0011001111001100001100111100110010100101010110101010010101011010,
64'b1001011010010110100101101001011011000011001111001100001100111100,
64'b0101101010100101101001010101101011110000111100001111000011110000,
64'b1001011001101001011010011001011011000011001111001100001100111100,
64'b0011001111001100001100111100110011111111000000001111111100000000,
64'b1100110011001100110011001100110010011001011001101001100101100110,
64'b1100110011001100110011001100110001010101101010100101010110101010,
64'b1001011010010110100101101001011001010101101010100101010110101010,
64'b1100001100111100110000110011110010100101010110101010010101011010,
64'b0011001111001100001100111100110011000011110000110011110000111100,
64'b0101101010100101101001010101101000111100001111000011110000111100,
64'b1100001100111100110000110011110001011010101001011010010101011010,
64'b1111000011110000111100001111000001101001011010011001011010010110,
64'b0000111100001111111100001111000001100110100110011001100101100110,
64'b1100001100111100110000110011110011110000000011110000111111110000,
64'b1100110000110011001100111100110011111111000000001111111100000000,
64'b1001011001101001011010011001011011110000000011110000111111110000,
64'b1010010110100101010110100101101011111111111111110000000000000000,
64'b1111000011110000111100001111000011000011110000110011110000111100,
64'b1111000011110000111100001111000000110011001100111100110011001100,
64'b1100001100111100110000110011110000110011001100111100110011001100,
64'b0000111111110000000011111111000000110011110011000011001111001100,
64'b0110100110010110011010011001011000001111000011111111000011110000,
64'b1111000011110000111100001111000001100110100110011001100101100110,
64'b0110100101101001100101101001011001011010010110100101101001011010,
64'b0101010101010101101010101010101001101001011010011001011010010110,
64'b0000000011111111111111110000000000000000111111111111111100000000,
64'b0110011001100110011001100110011001011010101001011010010101011010,
64'b1010010101011010101001010101101010011001100110010110011001100110,
64'b1010101001010101010101011010101011110000000011110000111111110000,
64'b0011001100110011110011001100110010011001100110010110011001100110,
64'b0110100101101001100101101001011010100101101001010101101001011010,
64'b0101101010100101101001010101101000110011001100111100110011001100,
64'b1111111111111111000000000000000001010101010101011010101010101010,
64'b0101010110101010010101011010101010010110100101101001011010010110,
64'b0101010101010101101010101010101001010101101010100101010110101010,
64'b0000111111110000000011111111000001101001011010011001011010010110,
64'b1010101001010101010101011010101010011001011001101001100101100110,
64'b0011001100110011110011001100110011000011001111001100001100111100,
64'b0101010110101010010101011010101001010101010101011010101010101010,
64'b1111000011110000111100001111000001100110100110011001100101100110,
64'b0110100101101001100101101001011010010110100101101001011010010110,
64'b1001100101100110100110010110011010101010010101010101010110101010,
64'b0110100101101001100101101001011010010110100101101001011010010110,
64'b0000000011111111111111110000000010011001011001101001100101100110,
64'b0011110000111100001111000011110001011010010110100101101001011010,
64'b0101010101010101101010101010101001100110011001100110011001100110,
64'b0011001111001100001100111100110001101001100101100110100110010110,
64'b0000111111110000000011111111000010011001100110010110011001100110,
64'b0101101010100101101001010101101011000011001111001100001100111100,
64'b0101101001011010010110100101101001101001011010011001011010010110,
64'b0000111100001111111100001111000011110000000011110000111111110000,
64'b1001100101100110100110010110011011001100110011001100110011001100,
64'b1001100101100110100110010110011001101001011010011001011010010110,
64'b0110011001100110011001100110011001101001100101100110100110010110,
64'b1100001100111100110000110011110000110011001100111100110011001100,
64'b1111000000001111000011111111000001101001100101100110100110010110,
64'b0011110000111100001111000011110011000011110000110011110000111100,
64'b1111111111111111000000000000000000110011110011000011001111001100,
64'b0011001100110011110011001100110000111100001111000011110000111100,
64'b0000111111110000000011111111000011000011001111001100001100111100,
64'b1010101001010101010101011010101000111100001111000011110000111100,
64'b1100110000110011001100111100110001011010101001011010010101011010,
64'b1001100101100110100110010110011011000011001111001100001100111100,
64'b1111111100000000111111110000000010101010010101010101010110101010,
64'b0110100101101001100101101001011001011010010110100101101001011010,
64'b1100001111000011001111000011110011000011001111001100001100111100,
64'b0011110000111100001111000011110010010110011010010110100110010110,
64'b1111000000001111000011111111000011110000111100001111000011110000,
64'b0000000011111111111111110000000010010110011010010110100110010110,
64'b1010010101011010101001010101101000001111111100000000111111110000,
64'b0000000000000000000000000000000010100101101001010101101001011010,
64'b0101101001011010010110100101101000001111111100000000111111110000,
64'b0101010110101010010101011010101000001111111100000000111111110000,
64'b0101101010100101101001010101101010100101010110101010010101011010,
64'b0101010101010101101010101010101011001100001100110011001111001100,
64'b0000000000000000000000000000000001011010101001011010010101011010,
64'b1010101010101010101010101010101000110011001100111100110011001100,
64'b1100001111000011001111000011110010011001011001101001100101100110,
64'b1100001100111100110000110011110011110000000011110000111111110000,
64'b0000000000000000000000000000000000111100110000111100001100111100,
64'b1010101010101010101010101010101001010101101010100101010110101010,
64'b0110011001100110011001100110011000111100110000111100001100111100,
64'b0000111111110000000011111111000010101010010101010101010110101010,
64'b0101101010100101101001010101101000110011110011000011001111001100,
64'b1100110000110011001100111100110010101010010101010101010110101010,
64'b1001100101100110100110010110011011111111000000001111111100000000,
64'b0000111100001111111100001111000001100110100110011001100101100110,
64'b1001011010010110100101101001011000001111000011111111000011110000,
64'b1100001111000011001111000011110001100110100110011001100101100110,
64'b1001100110011001011001100110011001011010010110100101101001011010,
64'b0000111100001111111100001111000001101001011010011001011010010110,
64'b0011110011000011110000110011110000000000111111111111111100000000,
64'b1010010101011010101001010101101001011010101001011010010101011010,
64'b0110011010011001100110010110011010011001100110010110011001100110,
64'b0000111100001111111100001111000011110000000011110000111111110000,
64'b0110100110010110011010011001011010011001100110010110011001100110,
64'b1001011010010110100101101001011010100101101001010101101001011010,
64'b0101101001011010010110100101101000110011001100111100110011001100,
64'b1100001100111100110000110011110010101010101010101010101010101010,
64'b1111111100000000111111110000000000000000111111111111111100000000,
64'b0110100110010110011010011001011010100101010110101010010101011010,
64'b0000111111110000000011111111000000000000000000000000000000000000,
64'b1001011010010110100101101001011011001100001100110011001111001100,
64'b0101010110101010010101011010101011000011110000110011110000111100,
64'b0101101010100101101001010101101000110011001100111100110011001100,
64'b0110011010011001100110010110011011000011110000110011110000111100,
64'b1100001111000011001111000011110000111100110000111100001100111100,
64'b0101010110101010010101011010101010011001011001101001100101100110,
64'b1001011001101001011010011001011011111111111111110000000000000000,
64'b1100001100111100110000110011110011000011110000110011110000111100,
64'b0011001111001100001100111100110010100101101001010101101001011010,
64'b0000111111110000000011111111000000110011110011000011001111001100,
64'b1001011001101001011010011001011010010110011010010110100110010110,
64'b1100110000110011001100111100110010010110011010010110100110010110,
64'b0110100110010110011010011001011001101001011010011001011010010110,
64'b1001011001101001011010011001011001011010010110100101101001011010,
64'b0011001111001100001100111100110010100101101001010101101001011010,
64'b1010101001010101010101011010101000111100001111000011110000111100,
64'b1100110000110011001100111100110000000000000000000000000000000000,
64'b0000111100001111111100001111000011110000111100001111000011110000,
64'b1010101010101010101010101010101001011010010110100101101001011010,
64'b0101010110101010010101011010101001101001011010011001011010010110,
64'b0000000000000000000000000000000011111111111111110000000000000000,
64'b1111000011110000111100001111000001100110100110011001100101100110,
64'b1010101010101010101010101010101000001111111100000000111111110000,
64'b0101010101010101101010101010101010010110011010010110100110010110,
64'b0101010101010101101010101010101010010110011010010110100110010110,
64'b1111111100000000111111110000000001101001100101100110100110010110,
64'b0110100110010110011010011001011010011001011001101001100101100110,
64'b1010010101011010101001010101101000110011110011000011001111001100,
64'b0101010101010101101010101010101010100101010110101010010101011010,
64'b0000000011111111111111110000000000000000000000000000000000000000,
64'b1111111111111111000000000000000011111111000000001111111100000000,
64'b0101010101010101101010101010101000110011110011000011001111001100,
64'b0101101001011010010110100101101011000011001111001100001100111100,
64'b0101101010100101101001010101101010101010101010101010101010101010,
64'b0000000011111111111111110000000001101001011010011001011010010110,
64'b1001100101100110100110010110011001010101101010100101010110101010,
64'b1100110011001100110011001100110000111100110000111100001100111100,
64'b0110011001100110011001100110011010010110011010010110100110010110,
64'b0101010101010101101010101010101010010110011010010110100110010110,
64'b0011110011000011110000110011110011000011110000110011110000111100,
64'b1100110000110011001100111100110000001111000011111111000011110000,
64'b1100110011001100110011001100110011001100001100110011001111001100,
64'b0101010101010101101010101010101000000000000000000000000000000000,
64'b1010101010101010101010101010101011111111111111110000000000000000,
64'b0110011001100110011001100110011000001111000011111111000011110000,
64'b1001100101100110100110010110011011110000000011110000111111110000,
64'b1100110000110011001100111100110011001100110011001100110011001100,
64'b0101010101010101101010101010101011000011001111001100001100111100,
64'b1001011010010110100101101001011001100110011001100110011001100110,
64'b1001100101100110100110010110011000110011001100111100110011001100,
64'b1100110011001100110011001100110001100110100110011001100101100110,
64'b1010010110100101010110100101101011111111000000001111111100000000,
64'b0000111111110000000011111111000011110000000011110000111111110000,
64'b1010010101011010101001010101101001010101010101011010101010101010,
64'b0011110000111100001111000011110011000011110000110011110000111100,
64'b0110100110010110011010011001011000001111111100000000111111110000,
64'b1100110000110011001100111100110010101010010101010101010110101010,
64'b0000111100001111111100001111000001100110100110011001100101100110,
64'b1010101010101010101010101010101011000011001111001100001100111100,
64'b0101010110101010010101011010101000000000111111111111111100000000,
64'b1001100110011001011001100110011000001111111100000000111111110000,
64'b0011110000111100001111000011110001101001100101100110100110010110,
64'b0000000011111111111111110000000011110000111100001111000011110000,
64'b0000000000000000000000000000000001101001011010011001011010010110,
64'b0101101010100101101001010101101001010101010101011010101010101010,
64'b1111111100000000111111110000000000000000111111111111111100000000,
64'b1100110011001100110011001100110001100110011001100110011001100110,
64'b0110100110010110011010011001011010100101010110101010010101011010,
64'b1001100110011001011001100110011010101010010101010101010110101010,
64'b1010010101011010101001010101101000110011001100111100110011001100,
64'b0110011010011001100110010110011001101001011010011001011010010110,
64'b0000111100001111111100001111000001011010101001011010010101011010,
64'b0110100110010110011010011001011011111111111111110000000000000000,
64'b1100001111000011001111000011110010101010010101010101010110101010,
64'b1111000011110000111100001111000011000011001111001100001100111100,
64'b1001011001101001011010011001011011111111000000001111111100000000,
64'b0101101001011010010110100101101011000011001111001100001100111100,
64'b1010010101011010101001010101101001100110011001100110011001100110,
64'b0000000000000000000000000000000001010101010101011010101010101010,
64'b1111000000001111000011111111000010010110100101101001011010010110,
64'b0101101010100101101001010101101011001100001100110011001111001100,
64'b1001100101100110100110010110011000110011001100111100110011001100,
64'b1100110011001100110011001100110001011010010110100101101001011010,
64'b1111000011110000111100001111000001101001100101100110100110010110,
64'b0011110011000011110000110011110001100110100110011001100101100110,
64'b1100110011001100110011001100110010101010101010101010101010101010,
64'b1111000000001111000011111111000010011001100110010110011001100110,
64'b0000000000000000000000000000000010100101010110101010010101011010,
64'b1001011001101001011010011001011001010101010101011010101010101010,
64'b1001100101100110100110010110011011110000000011110000111111110000,
64'b1100110000110011001100111100110000111100001111000011110000111100,
64'b0000000000000000000000000000000011001100110011001100110011001100,
64'b0000000011111111111111110000000001101001100101100110100110010110,
64'b0110011010011001100110010110011000001111000011111111000011110000,
64'b0110100101101001100101101001011001011010010110100101101001011010,
64'b1111000011110000111100001111000010011001011001101001100101100110,
64'b1111111100000000111111110000000000111100110000111100001100111100,
64'b1111000000001111000011111111000011000011110000110011110000111100,
64'b0101101001011010010110100101101001100110011001100110011001100110,
64'b0000000011111111111111110000000000111100001111000011110000111100,
64'b1010101010101010101010101010101010011001011001101001100101100110,
64'b0011110011000011110000110011110001100110011001100110011001100110,
64'b0110100101101001100101101001011010101010010101010101010110101010,
64'b0000111100001111111100001111000010100101010110101010010101011010,
64'b1010101010101010101010101010101011110000111100001111000011110000,
64'b1111111111111111000000000000000000111100110000111100001100111100,
64'b0110100101101001100101101001011011111111000000001111111100000000,
64'b0110100110010110011010011001011010011001011001101001100101100110,
64'b0101010110101010010101011010101011000011110000110011110000111100,
64'b1111111111111111000000000000000011110000000011110000111111110000,
64'b0000000011111111111111110000000010100101010110101010010101011010,
64'b1001100101100110100110010110011010010110100101101001011010010110,
64'b1111111111111111000000000000000000001111111100000000111111110000,
64'b0110011001100110011001100110011000111100001111000011110000111100,
64'b0101101010100101101001010101101010010110100101101001011010010110,
64'b0110100110010110011010011001011000110011001100111100110011001100,
64'b0101010110101010010101011010101001100110100110011001100101100110,
64'b0110011001100110011001100110011011111111000000001111111100000000,
64'b0000000000000000000000000000000011110000000011110000111111110000,
64'b0110100110010110011010011001011001010101010101011010101010101010,
64'b1001011001101001011010011001011011000011110000110011110000111100,
64'b0011001100110011110011001100110000001111111100000000111111110000,
64'b0000000000000000000000000000000010101010010101010101010110101010,
64'b0101010101010101101010101010101001100110100110011001100101100110,
64'b0110100101101001100101101001011011000011001111001100001100111100,
64'b0000000000000000000000000000000000000000111111111111111100000000,
64'b1001011010010110100101101001011000001111111100000000111111110000,
64'b0101101010100101101001010101101010100101010110101010010101011010,
64'b0110100101101001100101101001011011001100110011001100110011001100,
64'b0011001100110011110011001100110010101010101010101010101010101010,
64'b0110011001100110011001100110011001100110100110011001100101100110,
64'b1111111100000000111111110000000000001111000011111111000011110000,
64'b1111111111111111000000000000000000110011110011000011001111001100,
64'b1100110000110011001100111100110001010101010101011010101010101010,
64'b1111000011110000111100001111000010010110100101101001011010010110,
64'b1001100101100110100110010110011000000000111111111111111100000000,
64'b1100110011001100110011001100110001010101101010100101010110101010,
64'b0101101001011010010110100101101000000000000000000000000000000000,
64'b0101010110101010010101011010101000000000111111111111111100000000,
64'b0011110000111100001111000011110010011001011001101001100101100110,
64'b0011110000111100001111000011110011001100001100110011001111001100,
64'b0000000011111111111111110000000011110000111100001111000011110000,
64'b0110100101101001100101101001011011001100110011001100110011001100,
64'b1111000011110000111100001111000011000011110000110011110000111100,
64'b0000000011111111111111110000000001010101101010100101010110101010,
64'b1111111111111111000000000000000010100101101001010101101001011010,
64'b0110100110010110011010011001011011001100110011001100110011001100,
64'b1010010101011010101001010101101001101001100101100110100110010110,
64'b0101101010100101101001010101101011111111111111110000000000000000,
64'b0011110000111100001111000011110010011001100110010110011001100110,
64'b0110100110010110011010011001011000000000000000000000000000000000,
64'b0110011010011001100110010110011011111111111111110000000000000000,
64'b0011001111001100001100111100110010010110100101101001011010010110,
64'b1111111111111111000000000000000010100101101001010101101001011010,
64'b1001011010010110100101101001011001010101101010100101010110101010,
64'b0101101010100101101001010101101011110000111100001111000011110000,
64'b0011001111001100001100111100110000001111111100000000111111110000,
64'b0000000011111111111111110000000010011001100110010110011001100110,
64'b0101010101010101101010101010101000110011110011000011001111001100,
64'b0101101001011010010110100101101001011010010110100101101001011010,
64'b0011110011000011110000110011110000111100110000111100001100111100,
64'b0101010101010101101010101010101000000000000000000000000000000000,
64'b0110100110010110011010011001011010010110100101101001011010010110,
64'b0110011010011001100110010110011010101010101010101010101010101010,
64'b1001011001101001011010011001011000000000000000000000000000000000,
64'b0110011001100110011001100110011001101001100101100110100110010110,
64'b1010101010101010101010101010101010011001011001101001100101100110,
64'b0110100110010110011010011001011010011001100110010110011001100110,
64'b1100110000110011001100111100110011111111000000001111111100000000,
64'b1010010110100101010110100101101000000000111111111111111100000000,
64'b1111111111111111000000000000000000111100001111000011110000111100,
64'b0110011001100110011001100110011010100101101001010101101001011010,
64'b1001100101100110100110010110011000110011110011000011001111001100,
64'b1111000000001111000011111111000011110000000011110000111111110000,
64'b0110011001100110011001100110011010101010101010101010101010101010,
64'b1001011001101001011010011001011011000011001111001100001100111100,
64'b1100001111000011001111000011110011001100110011001100110011001100,
64'b1001011001101001011010011001011000000000000000000000000000000000,
64'b1001011010010110100101101001011011000011001111001100001100111100,
64'b0011110011000011110000110011110001101001011010011001011010010110,
64'b0101010110101010010101011010101000111100001111000011110000111100,
64'b0011110000111100001111000011110001010101010101011010101010101010,
64'b1111111100000000111111110000000011111111111111110000000000000000,
64'b0101010110101010010101011010101010100101010110101010010101011010,
64'b0110100101101001100101101001011000110011110011000011001111001100,
64'b0000111111110000000011111111000010100101101001010101101001011010,
64'b1111000000001111000011111111000000000000111111111111111100000000,
64'b0000111111110000000011111111000001100110011001100110011001100110,
64'b1111000000001111000011111111000011110000000011110000111111110000,
64'b1111111100000000111111110000000011110000111100001111000011110000,
64'b1100001111000011001111000011110000000000000000000000000000000000,
64'b0101010110101010010101011010101000001111111100000000111111110000,
64'b0000000000000000000000000000000001101001100101100110100110010110,
64'b1111000011110000111100001111000010100101010110101010010101011010,
64'b0011110011000011110000110011110011001100110011001100110011001100,
64'b1001100110011001011001100110011010101010101010101010101010101010,
64'b1100110000110011001100111100110001100110100110011001100101100110,
64'b0011110011000011110000110011110000001111000011111111000011110000,
64'b0110011001100110011001100110011000110011110011000011001111001100,
64'b1111000000001111000011111111000001010101010101011010101010101010,
64'b0011001100110011110011001100110010010110100101101001011010010110,
64'b1100110000110011001100111100110000000000111111111111111100000000,
64'b0000111100001111111100001111000001010101101010100101010110101010,
64'b0101101001011010010110100101101000000000000000000000000000000000,
64'b0101101001011010010110100101101011111111000000001111111100000000,
64'b1010101010101010101010101010101001100110011001100110011001100110,
64'b1111111100000000111111110000000010100101010110101010010101011010,
64'b1111000000001111000011111111000011000011110000110011110000111100,
64'b1001011010010110100101101001011010101010101010101010101010101010,
64'b1010010110100101010110100101101000111100110000111100001100111100,
64'b0101101010100101101001010101101010101010010101010101010110101010,
64'b1001011010010110100101101001011001101001100101100110100110010110,
64'b0000000011111111111111110000000000111100001111000011110000111100,
64'b0101101001011010010110100101101011110000111100001111000011110000,
64'b1010010110100101010110100101101000110011001100111100110011001100,
64'b0101010110101010010101011010101011000011110000110011110000111100,
64'b1001100101100110100110010110011001010101101010100101010110101010,
64'b0011001111001100001100111100110000111100001111000011110000111100,
64'b0011110011000011110000110011110011001100001100110011001111001100,
64'b1001011010010110100101101001011010100101010110101010010101011010,
64'b0011001111001100001100111100110000111100110000111100001100111100,
64'b0000111111110000000011111111000000000000000000000000000000000000,
64'b1100110011001100110011001100110000001111000011111111000011110000,
64'b1001100101100110100110010110011001100110011001100110011001100110,
64'b1010010110100101010110100101101001011010010110100101101001011010,
64'b0000111100001111111100001111000011111111000000001111111100000000,
64'b0000000000000000000000000000000001100110011001100110011001100110,
64'b1111111100000000111111110000000000111100001111000011110000111100,
64'b1100001111000011001111000011110011111111000000001111111100000000,
64'b1001011001101001011010011001011011001100001100110011001111001100,
64'b1100110011001100110011001100110000110011110011000011001111001100,
64'b1010101010101010101010101010101010100101101001010101101001011010,
64'b0000000011111111111111110000000001100110100110011001100101100110,
64'b0011110000111100001111000011110011110000000011110000111111110000,
64'b0110011010011001100110010110011010101010101010101010101010101010,
64'b0000111111110000000011111111000011111111000000001111111100000000,
64'b0011110000111100001111000011110010010110100101101001011010010110,
64'b1111111111111111000000000000000000110011110011000011001111001100,
64'b1010010101011010101001010101101011111111111111110000000000000000,
64'b0011001111001100001100111100110000111100001111000011110000111100,
64'b0011001100110011110011001100110000001111111100000000111111110000,
64'b0101010110101010010101011010101011111111111111110000000000000000,
64'b1100001111000011001111000011110000001111000011111111000011110000,
64'b0110011001100110011001100110011001011010010110100101101001011010,
64'b0110011001100110011001100110011010011001011001101001100101100110,
64'b1111111111111111000000000000000001101001011010011001011010010110,
64'b1010010101011010101001010101101010101010010101010101010110101010,
64'b1100001111000011001111000011110001100110011001100110011001100110,
64'b1010101001010101010101011010101011111111111111110000000000000000,
64'b0000111111110000000011111111000011000011001111001100001100111100,
64'b0000000000000000000000000000000000001111000011111111000011110000,
64'b0110011010011001100110010110011000000000000000000000000000000000,
64'b0000111100001111111100001111000010100101010110101010010101011010,
64'b1111000011110000111100001111000000000000111111111111111100000000,
64'b1001100110011001011001100110011000000000000000000000000000000000,
64'b0000111111110000000011111111000001010101101010100101010110101010,
64'b1001011010010110100101101001011010011001011001101001100101100110,
64'b0110011010011001100110010110011010011001011001101001100101100110,
64'b0110100101101001100101101001011010101010010101010101010110101010,
64'b0101010110101010010101011010101010101010101010101010101010101010,
64'b0110100110010110011010011001011011110000111100001111000011110000,
64'b0110011010011001100110010110011011111111000000001111111100000000,
64'b0101010110101010010101011010101010100101010110101010010101011010,
64'b1100110000110011001100111100110000110011001100111100110011001100,
64'b0011001100110011110011001100110001011010010110100101101001011010,
64'b1100110011001100110011001100110001010101010101011010101010101010,
64'b1001100101100110100110010110011000110011001100111100110011001100,
64'b0110011001100110011001100110011011110000111100001111000011110000,
64'b1111111111111111000000000000000001100110100110011001100101100110,
64'b1111111100000000111111110000000000000000000000000000000000000000,
64'b1001100101100110100110010110011001101001011010011001011010010110,
64'b0000000011111111111111110000000000110011001100111100110011001100,
64'b1010101010101010101010101010101001100110011001100110011001100110,
64'b0101101010100101101001010101101011111111000000001111111100000000,
64'b0011110011000011110000110011110011111111111111110000000000000000,
64'b0110011001100110011001100110011011001100001100110011001111001100,
64'b1100001100111100110000110011110011110000111100001111000011110000,
64'b1010101010101010101010101010101010011001011001101001100101100110,
64'b1100001100111100110000110011110011001100110011001100110011001100,
64'b0000111100001111111100001111000001011010010110100101101001011010,
64'b0110011001100110011001100110011001010101101010100101010110101010,
64'b0101010110101010010101011010101011000011110000110011110000111100,
64'b1001011010010110100101101001011010101010101010101010101010101010,
64'b1001100101100110100110010110011001101001100101100110100110010110,
64'b1001011010010110100101101001011001011010010110100101101001011010,
64'b0101010101010101101010101010101010010110100101101001011010010110,
64'b1010101001010101010101011010101011111111111111110000000000000000,
64'b1010010110100101010110100101101000000000000000000000000000000000,
64'b0110100101101001100101101001011010100101101001010101101001011010,
64'b0011110000111100001111000011110001010101101010100101010110101010,
64'b0011110000111100001111000011110011000011110000110011110000111100,
64'b0110100101101001100101101001011011110000111100001111000011110000,
64'b0011001111001100001100111100110000110011110011000011001111001100,
64'b1100110011001100110011001100110000110011001100111100110011001100,
64'b0110011010011001100110010110011000001111111100000000111111110000,
64'b1111111100000000111111110000000001100110011001100110011001100110,
64'b1100001111000011001111000011110010010110011010010110100110010110,
64'b1100001100111100110000110011110000110011110011000011001111001100,
64'b1100110011001100110011001100110011000011001111001100001100111100,
64'b1001100110011001011001100110011000000000000000000000000000000000,
64'b1001100101100110100110010110011010101010101010101010101010101010,
64'b0110100110010110011010011001011000110011110011000011001111001100,
64'b1010010101011010101001010101101010011001100110010110011001100110,
64'b0000111111110000000011111111000000001111111100000000111111110000,
64'b1100001100111100110000110011110001010101101010100101010110101010,
64'b1010010110100101010110100101101000001111000011111111000011110000,
64'b1111000011110000111100001111000011110000111100001111000011110000,
64'b1100001111000011001111000011110010101010010101010101010110101010,
64'b1010101010101010101010101010101000111100001111000011110000111100,
64'b0000111111110000000011111111000010010110011010010110100110010110,
64'b0101101010100101101001010101101010100101101001010101101001011010,
64'b1111000011110000111100001111000011110000000011110000111111110000,
64'b0011110000111100001111000011110000000000000000000000000000000000,
64'b0110100101101001100101101001011011001100110011001100110011001100,
64'b0011110011000011110000110011110000001111000011111111000011110000,
64'b1100110000110011001100111100110000111100001111000011110000111100,
64'b0000000011111111111111110000000010101010010101010101010110101010,
64'b1111000000001111000011111111000000110011001100111100110011001100,
64'b0011001111001100001100111100110011111111000000001111111100000000,
64'b0101010110101010010101011010101001010101101010100101010110101010,
64'b0000111111110000000011111111000000110011001100111100110011001100,
64'b0110011001100110011001100110011010100101010110101010010101011010,
64'b0000000011111111111111110000000000111100110000111100001100111100,
64'b1100110000110011001100111100110010011001011001101001100101100110,
64'b0101010110101010010101011010101010101010010101010101010110101010,
64'b0000111111110000000011111111000010101010101010101010101010101010,
64'b1100001100111100110000110011110011110000111100001111000011110000,
64'b0101101010100101101001010101101011111111000000001111111100000000,
64'b1010010110100101010110100101101010100101010110101010010101011010,
64'b0101010101010101101010101010101000110011001100111100110011001100,
64'b1010101001010101010101011010101001011010010110100101101001011010,
64'b1010010110100101010110100101101001010101010101011010101010101010,
64'b0011001100110011110011001100110000110011001100111100110011001100,
64'b0000000011111111111111110000000011110000111100001111000011110000,
64'b0011110000111100001111000011110010011001011001101001100101100110,
64'b0110011001100110011001100110011001100110100110011001100101100110,
64'b1111000000001111000011111111000010101010101010101010101010101010,
64'b1010010110100101010110100101101000111100001111000011110000111100,
64'b0011110011000011110000110011110001101001011010011001011010010110,
64'b1010101010101010101010101010101011110000111100001111000011110000,
64'b1100001100111100110000110011110001101001100101100110100110010110,
64'b1001100110011001011001100110011000111100110000111100001100111100,
64'b1100001111000011001111000011110000000000000000000000000000000000,
64'b0101010110101010010101011010101011001100001100110011001111001100,
64'b1100110011001100110011001100110010101010101010101010101010101010,
64'b1111111100000000111111110000000000001111111100000000111111110000,
64'b1001011010010110100101101001011010101010010101010101010110101010,
64'b1010101010101010101010101010101011001100110011001100110011001100,
64'b0101101001011010010110100101101001101001011010011001011010010110,
64'b1111000011110000111100001111000001100110011001100110011001100110,
64'b0011110011000011110000110011110000001111111100000000111111110000,
64'b0110011001100110011001100110011011000011001111001100001100111100,
64'b1100110011001100110011001100110001010101101010100101010110101010,
64'b0011001100110011110011001100110000111100110000111100001100111100,
64'b1010010110100101010110100101101011110000000011110000111111110000,
64'b0110011010011001100110010110011010101010101010101010101010101010,
64'b1100110000110011001100111100110000001111000011111111000011110000,
64'b0011110000111100001111000011110001100110011001100110011001100110,
64'b0000000011111111111111110000000000000000111111111111111100000000,
64'b0101010110101010010101011010101000110011001100111100110011001100,
64'b0110011001100110011001100110011001011010010110100101101001011010,
64'b1111111100000000111111110000000011000011001111001100001100111100,
64'b0000111100001111111100001111000010010110100101101001011010010110,
64'b0101010110101010010101011010101000000000111111111111111100000000,
64'b1010101001010101010101011010101011110000000011110000111111110000,
64'b0101101001011010010110100101101000110011001100111100110011001100,
64'b0011001111001100001100111100110011110000000011110000111111110000,
64'b0000000011111111111111110000000010101010010101010101010110101010,
64'b1010101010101010101010101010101001100110011001100110011001100110,
64'b1111000000001111000011111111000011111111000000001111111100000000,
64'b0110100110010110011010011001011010010110100101101001011010010110,
64'b0000000011111111111111110000000011111111111111110000000000000000,
64'b0000111100001111111100001111000001011010010110100101101001011010,
64'b1001011010010110100101101001011010011001011001101001100101100110,
64'b1111111111111111000000000000000001011010101001011010010101011010,
64'b1111111100000000111111110000000011000011001111001100001100111100,
64'b1001100110011001011001100110011011111111111111110000000000000000,
64'b0011001100110011110011001100110010101010010101010101010110101010,
64'b1001100101100110100110010110011001011010010110100101101001011010,
64'b0000111100001111111100001111000010101010010101010101010110101010,
64'b1111111111111111000000000000000010011001100110010110011001100110,
64'b0110011001100110011001100110011010010110100101101001011010010110,
64'b0000000011111111111111110000000011111111111111110000000000000000,
64'b1001011001101001011010011001011011000011001111001100001100111100,
64'b1111111111111111000000000000000000000000000000000000000000000000,
64'b0101010110101010010101011010101010011001011001101001100101100110,
64'b0110100110010110011010011001011000111100001111000011110000111100,
64'b0110011001100110011001100110011001100110100110011001100101100110,
64'b1010010101011010101001010101101001011010101001011010010101011010,
64'b1001100110011001011001100110011000000000000000000000000000000000,
64'b0110011010011001100110010110011010011001100110010110011001100110,
64'b1100001111000011001111000011110010011001011001101001100101100110,
64'b0011110000111100001111000011110000110011001100111100110011001100,
64'b0011001100110011110011001100110010010110100101101001011010010110,
64'b0101010101010101101010101010101001101001100101100110100110010110,
64'b1010101001010101010101011010101000000000000000000000000000000000,
64'b0101101010100101101001010101101001011010101001011010010101011010,
64'b0101010110101010010101011010101000000000000000000000000000000000,
64'b0000111100001111111100001111000011000011110000110011110000111100,
64'b0110100110010110011010011001011000001111111100000000111111110000,
64'b1111000011110000111100001111000001101001011010011001011010010110,
64'b0011110000111100001111000011110001100110100110011001100101100110,
64'b1001100110011001011001100110011010101010101010101010101010101010,
64'b0101010110101010010101011010101000111100001111000011110000111100,
64'b0000111111110000000011111111000001101001011010011001011010010110,
64'b0110011001100110011001100110011011110000111100001111000011110000,
64'b0110100101101001100101101001011001101001100101100110100110010110,
64'b1010010110100101010110100101101000111100110000111100001100111100,
64'b1100110000110011001100111100110000000000000000000000000000000000,
64'b1010101001010101010101011010101011001100001100110011001111001100,
64'b0110011010011001100110010110011010101010101010101010101010101010,
64'b0110100110010110011010011001011000001111111100000000111111110000,
64'b1100001100111100110000110011110001010101101010100101010110101010,
64'b1111111100000000111111110000000000001111111100000000111111110000,
64'b0000111111110000000011111111000010011001011001101001100101100110,
64'b0011110000111100001111000011110011000011110000110011110000111100,
64'b1001100110011001011001100110011000110011001100111100110011001100,
64'b0000000011111111111111110000000001101001100101100110100110010110,
64'b0011110000111100001111000011110010010110100101101001011010010110,
64'b1100001100111100110000110011110010100101010110101010010101011010,
64'b1001100101100110100110010110011000110011110011000011001111001100,
64'b1010010110100101010110100101101011111111000000001111111100000000,
64'b1001100110011001011001100110011011000011110000110011110000111100,
64'b0110100101101001100101101001011010011001011001101001100101100110,
64'b1001011001101001011010011001011010010110011010010110100110010110,
64'b0000111111110000000011111111000001100110011001100110011001100110,
64'b0011001100110011110011001100110001100110100110011001100101100110,
64'b1111000011110000111100001111000000110011110011000011001111001100,
64'b1010101001010101010101011010101010101010010101010101010110101010,
64'b0000000011111111111111110000000001100110100110011001100101100110,
64'b1111111111111111000000000000000000111100110000111100001100111100,
64'b0110011001100110011001100110011000000000000000000000000000000000,
64'b0110100110010110011010011001011001010101101010100101010110101010,
64'b0000000000000000000000000000000011001100110011001100110011001100,
64'b0110011001100110011001100110011010101010010101010101010110101010,
64'b0101101001011010010110100101101011000011001111001100001100111100,
64'b1001011010010110100101101001011010010110011010010110100110010110,
64'b0000000011111111111111110000000010101010010101010101010110101010,
64'b1111111100000000111111110000000000111100001111000011110000111100,
64'b1001011010010110100101101001011001101001011010011001011010010110,
64'b1010010110100101010110100101101010100101101001010101101001011010,
64'b1001011010010110100101101001011000110011001100111100110011001100,
64'b0110100110010110011010011001011001101001011010011001011010010110,
64'b0000000000000000000000000000000001011010101001011010010101011010,
64'b0101010110101010010101011010101010101010101010101010101010101010,
64'b1010010101011010101001010101101000110011001100111100110011001100,
64'b1100001111000011001111000011110011110000111100001111000011110000,
64'b0110100110010110011010011001011000110011001100111100110011001100,
64'b1111111100000000111111110000000001011010101001011010010101011010,
64'b0011110000111100001111000011110000111100110000111100001100111100,
64'b0110100101101001100101101001011010011001100110010110011001100110,
64'b0000000000000000000000000000000010100101010110101010010101011010,
64'b1100001100111100110000110011110011000011001111001100001100111100,
64'b0011001111001100001100111100110010011001011001101001100101100110,
64'b0110100110010110011010011001011001011010010110100101101001011010,
64'b0011110011000011110000110011110001101001100101100110100110010110,
64'b0000000000000000000000000000000001100110100110011001100101100110,
64'b0011001100110011110011001100110001100110011001100110011001100110,
64'b1100110000110011001100111100110011110000111100001111000011110000,
64'b0000111111110000000011111111000001010101101010100101010110101010,
64'b1001011001101001011010011001011011110000111100001111000011110000,
64'b1111111111111111000000000000000001100110100110011001100101100110,
64'b0000111111110000000011111111000001011010101001011010010101011010,
64'b1100001100111100110000110011110010010110100101101001011010010110,
64'b1010101010101010101010101010101010011001011001101001100101100110,
64'b1001011001101001011010011001011000111100110000111100001100111100,
64'b1111111100000000111111110000000000110011110011000011001111001100,
64'b1001100101100110100110010110011010010110011010010110100110010110,
64'b1100110011001100110011001100110000000000000000000000000000000000,
64'b0000000000000000000000000000000001101001011010011001011010010110,
64'b0011001111001100001100111100110001010101101010100101010110101010,
64'b0011110000111100001111000011110001100110100110011001100101100110,
64'b0110100110010110011010011001011011110000111100001111000011110000,
64'b0110100101101001100101101001011010101010101010101010101010101010,
64'b0110011001100110011001100110011000001111000011111111000011110000,
64'b0101010101010101101010101010101010011001100110010110011001100110,
64'b0110011010011001100110010110011011111111000000001111111100000000,
64'b0110011001100110011001100110011010010110100101101001011010010110,
64'b1111000000001111000011111111000011110000000011110000111111110000,
64'b1010010101011010101001010101101010100101101001010101101001011010,
64'b0110011001100110011001100110011000111100110000111100001100111100,
64'b1100110000110011001100111100110010101010101010101010101010101010,
64'b1010101010101010101010101010101011000011001111001100001100111100,
64'b1100110000110011001100111100110010011001100110010110011001100110,
64'b1001011001101001011010011001011011000011110000110011110000111100,
64'b1111111100000000111111110000000001010101101010100101010110101010,
64'b1001011010010110100101101001011011001100110011001100110011001100,
64'b0101101001011010010110100101101011111111000000001111111100000000,
64'b0011001111001100001100111100110010010110100101101001011010010110,
64'b1111111111111111000000000000000001010101010101011010101010101010,
64'b0011110000111100001111000011110011000011001111001100001100111100,
64'b0110011010011001100110010110011000000000111111111111111100000000,
64'b1001011010010110100101101001011010011001011001101001100101100110,
64'b1001100110011001011001100110011001011010101001011010010101011010,
64'b0011001111001100001100111100110001100110011001100110011001100110,
64'b1100110011001100110011001100110011110000000011110000111111110000,
64'b1100110000110011001100111100110000111100001111000011110000111100,
64'b0000111111110000000011111111000010100101010110101010010101011010,
64'b1001011010010110100101101001011010011001100110010110011001100110,
64'b1001011010010110100101101001011011110000111100001111000011110000,
64'b1111111100000000111111110000000011111111111111110000000000000000,
64'b1111000000001111000011111111000011000011001111001100001100111100,
64'b1001011010010110100101101001011011001100110011001100110011001100,
64'b0000111111110000000011111111000010100101010110101010010101011010,
64'b0110100101101001100101101001011011111111111111110000000000000000,
64'b0110100110010110011010011001011001101001011010011001011010010110,
64'b0011110000111100001111000011110011001100001100110011001111001100,
64'b1010010110100101010110100101101010010110100101101001011010010110,
64'b1111000011110000111100001111000000000000111111111111111100000000,
64'b0000111100001111111100001111000010100101010110101010010101011010,
64'b1010101001010101010101011010101011001100001100110011001111001100,
64'b1100001100111100110000110011110000111100001111000011110000111100,
64'b1100001100111100110000110011110001010101101010100101010110101010,
64'b1111111111111111000000000000000000000000000000000000000000000000,
64'b0000000011111111111111110000000001011010101001011010010101011010,
64'b0110100110010110011010011001011011110000111100001111000011110000,
64'b1111111100000000111111110000000000110011110011000011001111001100,
64'b1100001100111100110000110011110000000000000000000000000000000000,
64'b1001011001101001011010011001011001101001100101100110100110010110,
64'b0000111111110000000011111111000010100101101001010101101001011010,
64'b0011001111001100001100111100110001101001100101100110100110010110,
64'b0101010110101010010101011010101011111111111111110000000000000000,
64'b1111111100000000111111110000000001100110100110011001100101100110,
64'b1001100110011001011001100110011000001111000011111111000011110000,
64'b0101101010100101101001010101101010100101010110101010010101011010,
64'b1111000000001111000011111111000000110011001100111100110011001100,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0101010101010101101010101010101011001100001100110011001111001100,
64'b1001011001101001011010011001011001010101101010100101010110101010,
64'b0000000000000000000000000000000011110000111100001111000011110000,
64'b1111000000001111000011111111000010101010101010101010101010101010,
64'b0011110011000011110000110011110000111100110000111100001100111100,
64'b1010101001010101010101011010101000110011110011000011001111001100,
64'b0000111100001111111100001111000010010110011010010110100110010110,
64'b0011001100110011110011001100110000000000000000000000000000000000,
64'b1111111111111111000000000000000001101001011010011001011010010110,
64'b0011110000111100001111000011110001010101101010100101010110101010,
64'b0110011010011001100110010110011001100110100110011001100101100110,
64'b1010101001010101010101011010101011110000111100001111000011110000,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b1100110011001100110011001100110000001111000011111111000011110000,
64'b1001011001101001011010011001011010011001100110010110011001100110,
64'b1010101010101010101010101010101011111111000000001111111100000000,
64'b0101101010100101101001010101101010101010101010101010101010101010,
64'b0000111111110000000011111111000001011010010110100101101001011010,
64'b1010101010101010101010101010101000110011001100111100110011001100,
64'b1100110000110011001100111100110010010110100101101001011010010110,
64'b1001011001101001011010011001011000000000111111111111111100000000,
64'b1111000000001111000011111111000001101001100101100110100110010110,
64'b0011110000111100001111000011110011000011110000110011110000111100,
64'b0110100110010110011010011001011010011001011001101001100101100110,
64'b0000111100001111111100001111000010100101101001010101101001011010,
64'b0000111111110000000011111111000011110000111100001111000011110000,
64'b1111111111111111000000000000000001100110011001100110011001100110,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000001101001100101100110100110010110,
64'b1001011010010110100101101001011011001100110011001100110011001100,
64'b1010010110100101010110100101101000110011110011000011001111001100,
64'b0110011001100110011001100110011011110000111100001111000011110000,
64'b1100001100111100110000110011110001101001100101100110100110010110,
64'b0000000000000000000000000000000011111111111111110000000000000000,
64'b0101101001011010010110100101101010010110011010010110100110010110,
64'b1001100101100110100110010110011000001111111100000000111111110000,
64'b0101010101010101101010101010101001101001011010011001011010010110,
64'b1111000000001111000011111111000000110011110011000011001111001100,
64'b1010010110100101010110100101101001010101101010100101010110101010,
64'b1111111111111111000000000000000000111100001111000011110000111100,
64'b1010101010101010101010101010101000000000000000000000000000000000,
64'b0000000000000000000000000000000011000011001111001100001100111100,
64'b1001100110011001011001100110011011110000111100001111000011110000,
64'b0011110000111100001111000011110000001111000011111111000011110000,
64'b0011110000111100001111000011110011111111000000001111111100000000,
64'b0011110000111100001111000011110000111100110000111100001100111100,
64'b1001011001101001011010011001011000000000000000000000000000000000,
64'b1100001111000011001111000011110010010110011010010110100110010110,
64'b1111111111111111000000000000000010101010010101010101010110101010,
64'b1010010101011010101001010101101011000011001111001100001100111100,
64'b1010010101011010101001010101101010100101101001010101101001011010,
64'b1001011010010110100101101001011000110011001100111100110011001100,
64'b0101010101010101101010101010101000001111111100000000111111110000,
64'b0110011001100110011001100110011000000000000000000000000000000000,
64'b0000000000000000000000000000000000001111111100000000111111110000,
64'b0011110000111100001111000011110001010101101010100101010110101010,
64'b1010010101011010101001010101101011111111000000001111111100000000,
64'b0000111111110000000011111111000001010101010101011010101010101010,
64'b0000111111110000000011111111000011110000000011110000111111110000,
64'b0011110011000011110000110011110010101010101010101010101010101010,
64'b1010010101011010101001010101101000111100110000111100001100111100,
64'b1010101010101010101010101010101010011001100110010110011001100110,
64'b0110011010011001100110010110011001011010101001011010010101011010,
64'b1100110000110011001100111100110000110011110011000011001111001100,
64'b1100001100111100110000110011110001011010010110100101101001011010,
64'b1100110011001100110011001100110010101010010101010101010110101010,
64'b1001011010010110100101101001011000000000000000000000000000000000,
64'b0000000000000000000000000000000011111111000000001111111100000000,
64'b1111111111111111000000000000000000110011001100111100110011001100,
64'b1100001111000011001111000011110011111111111111110000000000000000,
64'b1010101001010101010101011010101011001100110011001100110011001100,
64'b1100110011001100110011001100110010101010010101010101010110101010,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b1001011010010110100101101001011011110000000011110000111111110000,
64'b1111000011110000111100001111000010010110100101101001011010010110,
64'b1010101001010101010101011010101001100110100110011001100101100110,
64'b1010101010101010101010101010101010100101101001010101101001011010,
64'b0101010101010101101010101010101000110011110011000011001111001100,
64'b0000111100001111111100001111000000110011001100111100110011001100,
64'b1100001100111100110000110011110010101010101010101010101010101010,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1111000000001111000011111111000001011010010110100101101001011010,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b0011001100110011110011001100110001011010010110100101101001011010,
64'b1001011001101001011010011001011000110011001100111100110011001100,
64'b1010101001010101010101011010101010010110100101101001011010010110,
64'b0011001100110011110011001100110000000000111111111111111100000000,
64'b1100001100111100110000110011110001101001100101100110100110010110,
64'b0101101010100101101001010101101011000011110000110011110000111100,
64'b0110100101101001100101101001011010011001011001101001100101100110,
64'b1100001100111100110000110011110010100101101001010101101001011010,
64'b1010101001010101010101011010101011110000111100001111000011110000,
64'b0101101010100101101001010101101001100110011001100110011001100110,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1010101001010101010101011010101011000011110000110011110000111100,
64'b0110011001100110011001100110011011000011001111001100001100111100,
64'b1111000011110000111100001111000010011001011001101001100101100110,
64'b1001011001101001011010011001011000111100110000111100001100111100,
64'b1001100110011001011001100110011011111111111111110000000000000000,
64'b0101101001011010010110100101101000001111111100000000111111110000,
64'b0101101010100101101001010101101010101010010101010101010110101010,
64'b1100110000110011001100111100110001100110011001100110011001100110,
64'b0110100110010110011010011001011001100110011001100110011001100110,
64'b0101101010100101101001010101101000111100001111000011110000111100,
64'b0011001100110011110011001100110010101010010101010101010110101010,
64'b0110011010011001100110010110011000111100001111000011110000111100,
64'b1010101010101010101010101010101000000000000000000000000000000000,
64'b1100001100111100110000110011110001010101010101011010101010101010,
64'b1001100101100110100110010110011001010101010101011010101010101010,
64'b0101010110101010010101011010101001101001011010011001011010010110,
64'b1111000011110000111100001111000000111100001111000011110000111100,
64'b0000000011111111111111110000000000111100110000111100001100111100,
64'b0110100101101001100101101001011001011010010110100101101001011010,
64'b1111000000001111000011111111000000001111000011111111000011110000,
64'b1100110000110011001100111100110011111111000000001111111100000000,
64'b1001100101100110100110010110011000110011001100111100110011001100,
64'b1100001111000011001111000011110000000000000000000000000000000000,
64'b1010010110100101010110100101101011001100110011001100110011001100,
64'b0110100101101001100101101001011010100101010110101010010101011010,
64'b0110011001100110011001100110011000000000000000000000000000000000,
64'b0000000000000000000000000000000011001100110011001100110011001100,
64'b1100110000110011001100111100110001100110011001100110011001100110,
64'b1001100110011001011001100110011001101001100101100110100110010110,
64'b0011001100110011110011001100110010100101010110101010010101011010,
64'b0110100110010110011010011001011011110000000011110000111111110000,
64'b1001100110011001011001100110011010011001011001101001100101100110,
64'b1001011001101001011010011001011011111111000000001111111100000000,
64'b1100110000110011001100111100110001010101010101011010101010101010,
64'b0110011001100110011001100110011011110000111100001111000011110000,
64'b0000000000000000000000000000000010101010101010101010101010101010,
64'b0110011010011001100110010110011011110000111100001111000011110000,
64'b0110100110010110011010011001011011001100001100110011001111001100,
64'b1001011010010110100101101001011000000000000000000000000000000000,
64'b0000000000000000000000000000000001011010010110100101101001011010,
64'b0000111100001111111100001111000000111100001111000011110000111100,
64'b1001011010010110100101101001011000111100110000111100001100111100,
64'b0101101001011010010110100101101011001100001100110011001111001100,
64'b1001011001101001011010011001011000000000111111111111111100000000,
64'b0011110000111100001111000011110001101001011010011001011010010110,
64'b1001011001101001011010011001011011111111111111110000000000000000,
64'b1010010110100101010110100101101011001100110011001100110011001100,
64'b1001011010010110100101101001011001010101101010100101010110101010,
64'b0000000000000000000000000000000011001100110011001100110011001100,
64'b1100001111000011001111000011110011111111000000001111111100000000,
64'b1001011001101001011010011001011000001111000011111111000011110000,
64'b1100001100111100110000110011110010101010101010101010101010101010,
64'b0101101010100101101001010101101011000011110000110011110000111100,
64'b1111000011110000111100001111000000000000000000000000000000000000,
64'b1100001100111100110000110011110001011010101001011010010101011010,
64'b1111111111111111000000000000000001101001100101100110100110010110,
64'b1010101010101010101010101010101011000011001111001100001100111100,
64'b0101010101010101101010101010101010011001100110010110011001100110,
64'b0000000011111111111111110000000010010110100101101001011010010110,
64'b1111000011110000111100001111000000110011110011000011001111001100,
64'b0110011010011001100110010110011000111100001111000011110000111100,
64'b0000111111110000000011111111000011111111000000001111111100000000,
64'b1111000000001111000011111111000000000000000000000000000000000000,
64'b1001011001101001011010011001011011111111000000001111111100000000,
64'b1010010101011010101001010101101001100110011001100110011001100110,
64'b1001011010010110100101101001011000001111111100000000111111110000,
64'b0101101001011010010110100101101010101010101010101010101010101010,
64'b0101101010100101101001010101101011001100001100110011001111001100,
64'b1100110000110011001100111100110010010110011010010110100110010110,
64'b1111000000001111000011111111000011110000000011110000111111110000,
64'b0011110011000011110000110011110000111100001111000011110000111100,
64'b0110100101101001100101101001011001101001100101100110100110010110,
64'b0011110000111100001111000011110000001111000011111111000011110000,
64'b1100110011001100110011001100110000001111111100000000111111110000,
64'b1010010110100101010110100101101011111111111111110000000000000000,
64'b1111111100000000111111110000000000000000000000000000000000000000,
64'b1001011001101001011010011001011011111111111111110000000000000000,
64'b1001100101100110100110010110011000111100001111000011110000111100,
64'b1001100110011001011001100110011010101010010101010101010110101010,
64'b0011110000111100001111000011110011001100110011001100110011001100,
64'b0110011010011001100110010110011000001111000011111111000011110000,
64'b0110100110010110011010011001011010010110011010010110100110010110,
64'b0011110000111100001111000011110010101010010101010101010110101010,
64'b1010101010101010101010101010101010100101010110101010010101011010,
64'b0101010110101010010101011010101000111100110000111100001100111100,
64'b1100110011001100110011001100110011111111000000001111111100000000,
64'b1111111111111111000000000000000010101010010101010101010110101010,
64'b0011110000111100001111000011110000000000000000000000000000000000,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b0011110011000011110000110011110000000000000000000000000000000000,
64'b1001011010010110100101101001011010100101010110101010010101011010,
64'b1001011010010110100101101001011010011001100110010110011001100110,
64'b1010010101011010101001010101101001011010010110100101101001011010,
64'b1100001111000011001111000011110011111111000000001111111100000000,
64'b1001011001101001011010011001011010010110011010010110100110010110,
64'b0000111111110000000011111111000010011001100110010110011001100110,
64'b1100110011001100110011001100110001100110100110011001100101100110,
64'b0011001100110011110011001100110011110000000011110000111111110000,
64'b1111000011110000111100001111000001010101010101011010101010101010,
64'b0000000000000000000000000000000000110011001100111100110011001100,
64'b1010010101011010101001010101101010101010101010101010101010101010,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b1111000000001111000011111111000000000000000000000000000000000000,
64'b0110100110010110011010011001011000110011110011000011001111001100,
64'b0110100110010110011010011001011010010110100101101001011010010110,
64'b1100110000110011001100111100110010011001011001101001100101100110,
64'b0000111111110000000011111111000011111111111111110000000000000000,
64'b1001011001101001011010011001011000111100110000111100001100111100,
64'b1010101001010101010101011010101010010110100101101001011010010110,
64'b1111000011110000111100001111000001101001011010011001011010010110,
64'b1111000011110000111100001111000010101010010101010101010110101010,
64'b0101010110101010010101011010101001100110011001100110011001100110,
64'b0000000000000000000000000000000001011010010110100101101001011010,
64'b1100110000110011001100111100110001100110011001100110011001100110,
64'b1111000011110000111100001111000011110000111100001111000011110000,
64'b0000000011111111111111110000000000000000000000000000000000000000,
64'b0110100110010110011010011001011011110000111100001111000011110000,
64'b0011110011000011110000110011110011000011001111001100001100111100,
64'b0000111100001111111100001111000011000011110000110011110000111100,
64'b1010101001010101010101011010101000000000000000000000000000000000,
64'b0011110011000011110000110011110001011010101001011010010101011010,
64'b1001100110011001011001100110011001101001100101100110100110010110,
64'b0101010110101010010101011010101011000011001111001100001100111100,
64'b1111111100000000111111110000000010011001100110010110011001100110,
64'b0011001100110011110011001100110010010110100101101001011010010110,
64'b0000000000000000000000000000000000110011110011000011001111001100,
64'b0000111100001111111100001111000000111100001111000011110000111100,
64'b0101010110101010010101011010101011111111000000001111111100000000,
64'b1111111111111111000000000000000000000000000000000000000000000000,
64'b0110100110010110011010011001011011111111000000001111111100000000,
64'b1010010101011010101001010101101000110011110011000011001111001100,
64'b0011001111001100001100111100110000000000000000000000000000000000,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b0000111111110000000011111111000010011001011001101001100101100110,
64'b1100110000110011001100111100110001010101101010100101010110101010,
64'b0000000011111111111111110000000011001100110011001100110011001100,
64'b1111111111111111000000000000000001010101010101011010101010101010,
64'b1001011010010110100101101001011010100101101001010101101001011010,
64'b0110011001100110011001100110011001100110100110011001100101100110,
64'b1111111111111111000000000000000000111100001111000011110000111100,
64'b0101010110101010010101011010101001010101010101011010101010101010,
64'b0000111111110000000011111111000011001100110011001100110011001100,
64'b1111111100000000111111110000000010101010101010101010101010101010,
64'b0110100101101001100101101001011010100101101001010101101001011010,
64'b0011110011000011110000110011110000000000000000000000000000000000,
64'b0101101001011010010110100101101000111100001111000011110000111100,
64'b0000111100001111111100001111000011000011110000110011110000111100,
64'b1100001100111100110000110011110000110011001100111100110011001100,
64'b0101010110101010010101011010101011110000111100001111000011110000,
64'b0101010101010101101010101010101011001100110011001100110011001100,
64'b1111111100000000111111110000000010011001011001101001100101100110,
64'b0101101001011010010110100101101001101001011010011001011010010110,
64'b1111111111111111000000000000000010100101010110101010010101011010,
64'b1100110000110011001100111100110011001100110011001100110011001100,
64'b0000111100001111111100001111000001011010010110100101101001011010,
64'b1111111100000000111111110000000011001100110011001100110011001100,
64'b0110011001100110011001100110011010011001011001101001100101100110,
64'b0110100101101001100101101001011010101010101010101010101010101010,
64'b1111111100000000111111110000000000001111111100000000111111110000,
64'b1111000011110000111100001111000000001111111100000000111111110000,
64'b1001011010010110100101101001011001011010010110100101101001011010,
64'b0011001111001100001100111100110001010101101010100101010110101010,
64'b0011001100110011110011001100110011110000111100001111000011110000,
64'b1100001111000011001111000011110011000011110000110011110000111100,
64'b0101010110101010010101011010101011000011001111001100001100111100,
64'b1111111111111111000000000000000001100110100110011001100101100110,
64'b1111000000001111000011111111000011110000111100001111000011110000,
64'b0101101001011010010110100101101000110011110011000011001111001100,
64'b0101010110101010010101011010101011110000111100001111000011110000,
64'b0011110000111100001111000011110001101001011010011001011010010110,
64'b1100001100111100110000110011110011001100110011001100110011001100,
64'b0101010101010101101010101010101000000000111111111111111100000000,
64'b1111111100000000111111110000000000000000111111111111111100000000,
64'b1100001100111100110000110011110000110011110011000011001111001100,
64'b0000111100001111111100001111000000110011001100111100110011001100,
64'b1111000011110000111100001111000011111111000000001111111100000000,
64'b1010010101011010101001010101101000001111111100000000111111110000,
64'b1001100110011001011001100110011001011010101001011010010101011010,
64'b0000000000000000000000000000000011000011110000110011110000111100,
64'b1010101001010101010101011010101001010101101010100101010110101010,
64'b1001100101100110100110010110011000001111000011111111000011110000,
64'b1100110011001100110011001100110011111111000000001111111100000000,
64'b1010101010101010101010101010101001101001100101100110100110010110,
64'b1100001111000011001111000011110001011010010110100101101001011010,
64'b1010101010101010101010101010101011111111111111110000000000000000,
64'b0101101010100101101001010101101001010101010101011010101010101010,
64'b0011110000111100001111000011110010100101101001010101101001011010,
64'b1111111111111111000000000000000011110000111100001111000011110000,
64'b1010101001010101010101011010101001010101010101011010101010101010,
64'b0101101010100101101001010101101000000000111111111111111100000000,
64'b0101101001011010010110100101101011001100001100110011001111001100,
64'b0101010101010101101010101010101010100101010110101010010101011010,
64'b0110011010011001100110010110011010011001100110010110011001100110,
64'b0110011010011001100110010110011011111111000000001111111100000000,
64'b0000111111110000000011111111000010101010101010101010101010101010,
64'b0110100110010110011010011001011000111100110000111100001100111100,
64'b0011110000111100001111000011110000110011110011000011001111001100,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1100001111000011001111000011110001100110011001100110011001100110,
64'b0110100101101001100101101001011010011001011001101001100101100110,
64'b0000000011111111111111110000000001010101101010100101010110101010,
64'b0110011001100110011001100110011011001100110011001100110011001100,
64'b1111000000001111000011111111000001010101010101011010101010101010,
64'b1111111100000000111111110000000010100101101001010101101001011010,
64'b0011001100110011110011001100110001100110100110011001100101100110,
64'b0011110011000011110000110011110000111100001111000011110000111100,
64'b0110011010011001100110010110011001010101010101011010101010101010,
64'b1010101010101010101010101010101011001100110011001100110011001100,
64'b0011110011000011110000110011110001010101010101011010101010101010,
64'b0000111111110000000011111111000010010110011010010110100110010110,
64'b0000000000000000000000000000000001100110011001100110011001100110,
64'b0000111111110000000011111111000000110011110011000011001111001100,
64'b0110100110010110011010011001011000001111111100000000111111110000,
64'b0101010101010101101010101010101000110011110011000011001111001100,
64'b1001011010010110100101101001011000001111000011111111000011110000,
64'b0000000011111111111111110000000001011010010110100101101001011010,
64'b0101010101010101101010101010101011111111000000001111111100000000,
64'b1111000011110000111100001111000010010110100101101001011010010110,
64'b0101101010100101101001010101101011110000111100001111000011110000,
64'b0110100101101001100101101001011011000011001111001100001100111100,
64'b0110011001100110011001100110011010100101010110101010010101011010,
64'b0101010101010101101010101010101001101001100101100110100110010110,
64'b1001100110011001011001100110011010100101101001010101101001011010,
64'b0110011001100110011001100110011011110000111100001111000011110000,
64'b0000111100001111111100001111000000000000111111111111111100000000,
64'b1111000011110000111100001111000011001100110011001100110011001100,
64'b1100110000110011001100111100110000001111111100000000111111110000,
64'b1001011001101001011010011001011000000000111111111111111100000000,
64'b0110100101101001100101101001011000001111111100000000111111110000,
64'b0000000000000000000000000000000010011001100110010110011001100110,
64'b1010101001010101010101011010101000111100110000111100001100111100,
64'b1001100110011001011001100110011010101010101010101010101010101010,
64'b0110011001100110011001100110011011111111111111110000000000000000,
64'b0110100110010110011010011001011011001100110011001100110011001100,
64'b0110100110010110011010011001011000111100110000111100001100111100,
64'b1010010101011010101001010101101000110011110011000011001111001100,
64'b1111000011110000111100001111000001010101101010100101010110101010,
64'b1111000011110000111100001111000011111111111111110000000000000000,
64'b1001100110011001011001100110011001011010010110100101101001011010,
64'b0000111111110000000011111111000000000000111111111111111100000000,
64'b0110100110010110011010011001011011111111111111110000000000000000,
64'b1111111100000000111111110000000010101010010101010101010110101010,
64'b1100110011001100110011001100110000111100001111000011110000111100,
64'b1100110011001100110011001100110001011010101001011010010101011010,
64'b1100001100111100110000110011110001100110011001100110011001100110,
64'b1001100101100110100110010110011000000000000000000000000000000000,
64'b0011110000111100001111000011110001011010010110100101101001011010,
64'b0011110011000011110000110011110011110000000011110000111111110000,
64'b1100110000110011001100111100110010100101101001010101101001011010,
64'b1111111100000000111111110000000000110011001100111100110011001100,
64'b1111111100000000111111110000000000000000000000000000000000000000,
64'b0011110000111100001111000011110010011001011001101001100101100110,
64'b1010101001010101010101011010101011111111111111110000000000000000,
64'b0011110011000011110000110011110010101010101010101010101010101010,
64'b1111111111111111000000000000000010011001100110010110011001100110,
64'b1111000011110000111100001111000010100101010110101010010101011010,
64'b1111000011110000111100001111000011001100001100110011001111001100,
64'b1111000000001111000011111111000010010110100101101001011010010110,
64'b1100001111000011001111000011110000000000000000000000000000000000,
64'b0000111111110000000011111111000000110011110011000011001111001100,
64'b1111111111111111000000000000000010100101101001010101101001011010,
64'b1001011001101001011010011001011010101010101010101010101010101010,
64'b0011001100110011110011001100110000111100001111000011110000111100,
64'b1111000000001111000011111111000010100101010110101010010101011010,
64'b1100001111000011001111000011110000001111111100000000111111110000,
64'b0011001111001100001100111100110000000000111111111111111100000000,
64'b1010010101011010101001010101101010011001100110010110011001100110,
64'b0011110000111100001111000011110010101010101010101010101010101010,
64'b0011001111001100001100111100110000000000111111111111111100000000,
64'b0000000011111111111111110000000011110000111100001111000011110000,
64'b0101010101010101101010101010101000111100001111000011110000111100,
64'b1010101010101010101010101010101000001111111100000000111111110000,
64'b1010101010101010101010101010101000001111111100000000111111110000,
64'b0000111111110000000011111111000000110011110011000011001111001100,
64'b1010010110100101010110100101101001100110011001100110011001100110,
64'b0011110000111100001111000011110000001111111100000000111111110000,
64'b1010010110100101010110100101101011001100001100110011001111001100,
64'b0110100101101001100101101001011000000000111111111111111100000000,
64'b1010010101011010101001010101101011111111111111110000000000000000,
64'b0011001111001100001100111100110010010110100101101001011010010110,
64'b1001100101100110100110010110011001100110011001100110011001100110,
64'b0110100101101001100101101001011011111111111111110000000000000000,
64'b0000000000000000000000000000000001010101101010100101010110101010,
64'b0011001111001100001100111100110000001111111100000000111111110000,
64'b0110100110010110011010011001011000000000111111111111111100000000,
64'b0011001111001100001100111100110011111111000000001111111100000000,
64'b0000111100001111111100001111000000001111000011111111000011110000,
64'b0000000000000000000000000000000000111100001111000011110000111100,
64'b1100001100111100110000110011110000000000111111111111111100000000,
64'b0011110000111100001111000011110000001111000011111111000011110000,
64'b1010010110100101010110100101101001010101010101011010101010101010,
64'b0110011001100110011001100110011010101010101010101010101010101010,
64'b1111000011110000111100001111000001101001100101100110100110010110,
64'b0101010101010101101010101010101000111100001111000011110000111100,
64'b1010010101011010101001010101101000000000000000000000000000000000,
64'b0101010101010101101010101010101010011001100110010110011001100110,
64'b0101101010100101101001010101101000000000111111111111111100000000,
64'b0011001100110011110011001100110011111111111111110000000000000000,
64'b0000111111110000000011111111000010101010101010101010101010101010,
64'b1111111100000000111111110000000001010101101010100101010110101010,
64'b1010101010101010101010101010101010100101010110101010010101011010,
64'b1111000000001111000011111111000011111111111111110000000000000000,
64'b0000111111110000000011111111000001010101101010100101010110101010,
64'b0011001111001100001100111100110001100110011001100110011001100110,
64'b1001011010010110100101101001011001100110011001100110011001100110,
64'b1111111100000000111111110000000000111100110000111100001100111100,
64'b1100110011001100110011001100110000001111111100000000111111110000,
64'b0110011010011001100110010110011000000000000000000000000000000000,
64'b1100110011001100110011001100110000111100001111000011110000111100,
64'b0110011010011001100110010110011001010101010101011010101010101010,
64'b0101101001011010010110100101101010101010101010101010101010101010,
64'b0101010110101010010101011010101001100110011001100110011001100110,
64'b0101010101010101101010101010101010011001100110010110011001100110,
64'b1100110011001100110011001100110011001100001100110011001111001100,
64'b0000000011111111111111110000000000000000000000000000000000000000,
64'b1010101001010101010101011010101010011001100110010110011001100110,
64'b0000111100001111111100001111000000111100001111000011110000111100,
64'b1100001100111100110000110011110000111100001111000011110000111100,
64'b1111111111111111000000000000000011110000000011110000111111110000,
64'b1111000011110000111100001111000010101010010101010101010110101010,
64'b1100001111000011001111000011110000000000000000000000000000000000,
64'b0101101001011010010110100101101000001111111100000000111111110000,
64'b1100001111000011001111000011110011001100110011001100110011001100,
64'b1001100101100110100110010110011001100110011001100110011001100110,
64'b1100110011001100110011001100110000111100001111000011110000111100,
64'b0110011001100110011001100110011000111100001111000011110000111100,
64'b0101101001011010010110100101101010100101101001010101101001011010,
64'b1111111111111111000000000000000010101010101010101010101010101010,
64'b1001100110011001011001100110011000111100001111000011110000111100,
64'b0101010110101010010101011010101010100101010110101010010101011010,
64'b0101101010100101101001010101101000001111111100000000111111110000,
64'b0000000000000000000000000000000000000000111111111111111100000000,
64'b0101010110101010010101011010101010011001100110010110011001100110,
64'b0000111111110000000011111111000010101010101010101010101010101010,
64'b1001100101100110100110010110011000000000111111111111111100000000,
64'b0000111111110000000011111111000011110000111100001111000011110000,
64'b0110100101101001100101101001011000111100001111000011110000111100,
64'b1111000011110000111100001111000000001111111100000000111111110000,
64'b0101010101010101101010101010101001011010101001011010010101011010,
64'b1010101010101010101010101010101000000000111111111111111100000000,
64'b1100001100111100110000110011110000001111000011111111000011110000,
64'b1001011010010110100101101001011001011010101001011010010101011010,
64'b0011110000111100001111000011110000111100001111000011110000111100,
64'b1010101010101010101010101010101011110000000011110000111111110000,
64'b0000111111110000000011111111000010011001011001101001100101100110,
64'b0000111100001111111100001111000010101010010101010101010110101010,
64'b1100110000110011001100111100110011001100110011001100110011001100,
64'b1111000000001111000011111111000000110011110011000011001111001100,
64'b1111000000001111000011111111000010100101101001010101101001011010,
64'b1100001100111100110000110011110011110000111100001111000011110000,
64'b1001100101100110100110010110011010010110100101101001011010010110,
64'b0011001100110011110011001100110011001100001100110011001111001100,
64'b1100110011001100110011001100110001010101010101011010101010101010,
64'b0011001100110011110011001100110001010101101010100101010110101010,
64'b0101010110101010010101011010101001100110100110011001100101100110,
64'b0011001111001100001100111100110010100101010110101010010101011010,
64'b0110011001100110011001100110011000000000111111111111111100000000,
64'b0000111100001111111100001111000001101001011010011001011010010110,
64'b1111000000001111000011111111000000110011001100111100110011001100,
64'b0110100110010110011010011001011001011010010110100101101001011010,
64'b0101101001011010010110100101101000001111000011111111000011110000,
64'b0101101001011010010110100101101000110011110011000011001111001100,
64'b1001100110011001011001100110011001010101101010100101010110101010,
64'b1010010101011010101001010101101011000011001111001100001100111100,
64'b0000111100001111111100001111000000001111000011111111000011110000,
64'b1111000011110000111100001111000001100110011001100110011001100110,
64'b0011001111001100001100111100110010011001100110010110011001100110,
64'b0000111100001111111100001111000011000011110000110011110000111100,
64'b0011001100110011110011001100110001100110100110011001100101100110,
64'b1001011010010110100101101001011011111111111111110000000000000000,
64'b1111000011110000111100001111000001101001100101100110100110010110,
64'b1010010101011010101001010101101001011010010110100101101001011010,
64'b0101101001011010010110100101101010011001011001101001100101100110,
64'b1100001111000011001111000011110011111111000000001111111100000000,
64'b1100001111000011001111000011110010100101101001010101101001011010,
64'b1111111100000000111111110000000000110011001100111100110011001100,
64'b0000000000000000000000000000000000001111111100000000111111110000,
64'b0101010110101010010101011010101011111111000000001111111100000000,
64'b0101010110101010010101011010101010010110100101101001011010010110,
64'b0000111100001111111100001111000000111100001111000011110000111100,
64'b1111111100000000111111110000000010100101010110101010010101011010,
64'b0101101001011010010110100101101001101001011010011001011010010110,
64'b0110100110010110011010011001011010101010101010101010101010101010,
64'b1111111100000000111111110000000010010110011010010110100110010110,
64'b1100110000110011001100111100110000110011110011000011001111001100,
64'b0011001111001100001100111100110011000011110000110011110000111100,
64'b0000111111110000000011111111000011111111111111110000000000000000,
64'b1010010101011010101001010101101000110011110011000011001111001100,
64'b0101010101010101101010101010101001011010010110100101101001011010,
64'b0000000000000000000000000000000001010101101010100101010110101010,
64'b0110011001100110011001100110011001010101010101011010101010101010,
64'b1001100110011001011001100110011011000011001111001100001100111100,
64'b0011110000111100001111000011110000001111111100000000111111110000,
64'b1100001111000011001111000011110011001100001100110011001111001100,
64'b0000111111110000000011111111000011000011001111001100001100111100,
64'b1001011001101001011010011001011001100110011001100110011001100110,
64'b1111000000001111000011111111000000111100110000111100001100111100,
64'b0000000000000000000000000000000010100101101001010101101001011010,
64'b0110100110010110011010011001011000001111111100000000111111110000,
64'b1111000011110000111100001111000010101010101010101010101010101010,
64'b0011110000111100001111000011110010100101101001010101101001011010,
64'b0000111111110000000011111111000000110011110011000011001111001100,
64'b0011001111001100001100111100110011001100110011001100110011001100,
64'b1100001111000011001111000011110011001100110011001100110011001100,
64'b1001011010010110100101101001011001011010101001011010010101011010,
64'b0110011001100110011001100110011000000000111111111111111100000000,
64'b1001100101100110100110010110011000001111000011111111000011110000,
64'b1001011001101001011010011001011001011010101001011010010101011010,
64'b1001011001101001011010011001011000111100001111000011110000111100,
64'b1010010110100101010110100101101011110000000011110000111111110000,
64'b1010010110100101010110100101101010011001011001101001100101100110,
64'b1111000011110000111100001111000010101010010101010101010110101010,
64'b0000111100001111111100001111000011001100110011001100110011001100,
64'b1111111111111111000000000000000000110011110011000011001111001100,
64'b1100001111000011001111000011110010100101101001010101101001011010,
64'b0110100110010110011010011001011011110000111100001111000011110000,
64'b0000111111110000000011111111000010100101101001010101101001011010,
64'b0110100110010110011010011001011001100110100110011001100101100110,
64'b0011110000111100001111000011110010010110011010010110100110010110,
64'b1100001111000011001111000011110011000011001111001100001100111100,
64'b0011110011000011110000110011110001011010101001011010010101011010,
64'b1001011001101001011010011001011000001111111100000000111111110000,
64'b1001100101100110100110010110011000001111000011111111000011110000,
64'b1001100101100110100110010110011001100110011001100110011001100110,
64'b0101010110101010010101011010101011111111000000001111111100000000,
64'b1111111100000000111111110000000010101010010101010101010110101010,
64'b1010101010101010101010101010101011111111000000001111111100000000,
64'b1010010101011010101001010101101011110000111100001111000011110000,
64'b0110100110010110011010011001011011001100110011001100110011001100,
64'b0101010110101010010101011010101011001100001100110011001111001100,
64'b1001011001101001011010011001011011000011110000110011110000111100,
64'b1100110011001100110011001100110001010101010101011010101010101010,
64'b1001100101100110100110010110011011001100001100110011001111001100,
64'b0110011010011001100110010110011011110000000011110000111111110000,
64'b0011110011000011110000110011110000000000111111111111111100000000,
64'b0110011010011001100110010110011011110000111100001111000011110000,
64'b1100110011001100110011001100110010011001100110010110011001100110,
64'b1111111100000000111111110000000000110011110011000011001111001100,
64'b0000111111110000000011111111000011000011001111001100001100111100,
64'b0011110011000011110000110011110010100101010110101010010101011010,
64'b0000111100001111111100001111000000111100001111000011110000111100,
64'b0101101001011010010110100101101001101001100101100110100110010110,
64'b1100110011001100110011001100110000001111000011111111000011110000,
64'b1001011001101001011010011001011010100101010110101010010101011010,
64'b1001100101100110100110010110011001100110011001100110011001100110,
64'b0101010101010101101010101010101010100101101001010101101001011010,
64'b1111111111111111000000000000000010101010010101010101010110101010,
64'b1111000000001111000011111111000001010101010101011010101010101010,
64'b0110011010011001100110010110011001010101101010100101010110101010,
64'b0101010101010101101010101010101000111100001111000011110000111100,
64'b0011001111001100001100111100110010100101101001010101101001011010,
64'b1111000011110000111100001111000011110000000011110000111111110000,
64'b0000000000000000000000000000000011001100001100110011001111001100,
64'b1001011010010110100101101001011000001111111100000000111111110000,
64'b0000000000000000000000000000000011000011001111001100001100111100,
64'b1111000011110000111100001111000011111111000000001111111100000000,
64'b0011110011000011110000110011110001100110100110011001100101100110,
64'b0110100101101001100101101001011000111100001111000011110000111100,
64'b1100110011001100110011001100110000110011110011000011001111001100,
64'b1010101010101010101010101010101010011001100110010110011001100110,
64'b1010101001010101010101011010101001100110011001100110011001100110,
64'b0110100101101001100101101001011010011001100110010110011001100110,
64'b0110011001100110011001100110011000001111111100000000111111110000,
64'b1010010110100101010110100101101000110011110011000011001111001100,
64'b1111111100000000111111110000000010101010010101010101010110101010,
64'b0000000000000000000000000000000010100101101001010101101001011010,
64'b1100001100111100110000110011110010101010010101010101010110101010,
64'b0000000000000000000000000000000000001111111100000000111111110000,
64'b0000000011111111111111110000000000000000000000000000000000000000,
64'b0101101010100101101001010101101001101001011010011001011010010110,
64'b1010101010101010101010101010101001100110011001100110011001100110,
64'b1100110011001100110011001100110010011001100110010110011001100110,
64'b1111000011110000111100001111000000000000000000000000000000000000,
64'b1001100110011001011001100110011000111100001111000011110000111100,
64'b0110011001100110011001100110011000110011110011000011001111001100,
64'b1001100110011001011001100110011010100101010110101010010101011010,
64'b1111111111111111000000000000000011000011001111001100001100111100,
64'b1010010101011010101001010101101011000011001111001100001100111100,
64'b1111000000001111000011111111000001101001011010011001011010010110,
64'b0011001100110011110011001100110001011010101001011010010101011010,
64'b1001100101100110100110010110011011001100110011001100110011001100,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b1100110000110011001100111100110011000011001111001100001100111100,
64'b1010010101011010101001010101101010010110100101101001011010010110,
64'b0110011001100110011001100110011000111100001111000011110000111100,
64'b1100001100111100110000110011110010101010101010101010101010101010,
64'b1001011010010110100101101001011000001111111100000000111111110000,
64'b1001100101100110100110010110011000001111000011111111000011110000,
64'b0011001100110011110011001100110011001100001100110011001111001100,
64'b0110011010011001100110010110011011110000000011110000111111110000,
64'b1001011010010110100101101001011011110000000011110000111111110000,
64'b1111000011110000111100001111000011000011001111001100001100111100,
64'b1001100101100110100110010110011001100110100110011001100101100110,
64'b0000111111110000000011111111000001011010010110100101101001011010,
64'b0011001100110011110011001100110001100110011001100110011001100110,
64'b1010010110100101010110100101101011110000000011110000111111110000,
64'b1010010110100101010110100101101011000011001111001100001100111100,
64'b1010101010101010101010101010101000001111111100000000111111110000,
64'b1100110000110011001100111100110011001100110011001100110011001100,
64'b0110100110010110011010011001011000000000111111111111111100000000,
64'b1100110000110011001100111100110011111111000000001111111100000000,
64'b1111111111111111000000000000000010100101101001010101101001011010,
64'b1010010101011010101001010101101010101010010101010101010110101010,
64'b1001100110011001011001100110011010101010010101010101010110101010,
64'b0000111100001111111100001111000001011010101001011010010101011010,
64'b0000000011111111111111110000000011000011110000110011110000111100,
64'b0110011001100110011001100110011010011001011001101001100101100110,
64'b0101101001011010010110100101101000111100001111000011110000111100,
64'b1001100101100110100110010110011000000000111111111111111100000000,
64'b1001100101100110100110010110011001011010101001011010010101011010,
64'b0110011001100110011001100110011000000000111111111111111100000000,
64'b0000111100001111111100001111000011110000111100001111000011110000,
64'b1001011001101001011010011001011011111111111111110000000000000000,
64'b0000111100001111111100001111000001010101010101011010101010101010,
64'b1010101010101010101010101010101000110011110011000011001111001100,
64'b0110011010011001100110010110011010011001100110010110011001100110,
64'b0011110000111100001111000011110010011001100110010110011001100110,
64'b0101010110101010010101011010101001100110100110011001100101100110,
64'b0101010101010101101010101010101010100101010110101010010101011010,
64'b1001011010010110100101101001011010010110100101101001011010010110,
64'b1001100101100110100110010110011000001111111100000000111111110000,
64'b1100001111000011001111000011110011111111111111110000000000000000,
64'b1100001111000011001111000011110001100110100110011001100101100110,
64'b0011110000111100001111000011110001010101010101011010101010101010,
64'b1111111100000000111111110000000001010101101010100101010110101010,
64'b1001011001101001011010011001011000000000000000000000000000000000,
64'b0101010110101010010101011010101001100110011001100110011001100110,
64'b0110011001100110011001100110011010100101101001010101101001011010,
64'b1100001111000011001111000011110000111100001111000011110000111100,
64'b1010010101011010101001010101101010010110100101101001011010010110,
64'b0011001100110011110011001100110001101001011010011001011010010110,
64'b1100110011001100110011001100110001100110100110011001100101100110,
64'b0110100110010110011010011001011011000011001111001100001100111100,
64'b1100001111000011001111000011110000000000111111111111111100000000,
64'b0000111111110000000011111111000000000000000000000000000000000000,
64'b1010010101011010101001010101101001101001011010011001011010010110,
64'b1010010101011010101001010101101001100110011001100110011001100110,
64'b1111111111111111000000000000000010011001100110010110011001100110,
64'b0011110011000011110000110011110000000000000000000000000000000000,
64'b1001100110011001011001100110011000111100001111000011110000111100,
64'b0011110000111100001111000011110000110011110011000011001111001100,
64'b0000111111110000000011111111000010100101010110101010010101011010,
64'b0110011010011001100110010110011011000011001111001100001100111100,
64'b1111000011110000111100001111000011000011001111001100001100111100,
64'b0101101001011010010110100101101001101001011010011001011010010110,
64'b1100001100111100110000110011110010100101010110101010010101011010,
64'b1001100101100110100110010110011011111111000000001111111100000000,
64'b1111111100000000111111110000000001010101101010100101010110101010,
64'b1100110011001100110011001100110000000000000000000000000000000000,
64'b0000000011111111111111110000000010101010101010101010101010101010,
64'b1010101010101010101010101010101001011010010110100101101001011010,
64'b1001011010010110100101101001011011111111111111110000000000000000,
64'b0101101010100101101001010101101010010110011010010110100110010110,
64'b1111000011110000111100001111000001101001011010011001011010010110,
64'b1100110000110011001100111100110011111111000000001111111100000000,
64'b1010010101011010101001010101101000111100110000111100001100111100,
64'b1001100110011001011001100110011010011001100110010110011001100110,
64'b0000111111110000000011111111000011001100110011001100110011001100,
64'b0110100110010110011010011001011000110011110011000011001111001100,
64'b1111000000001111000011111111000011111111111111110000000000000000,
64'b0000000011111111111111110000000000110011001100111100110011001100,
64'b0011110000111100001111000011110000000000000000000000000000000000,
64'b1111111100000000111111110000000011001100110011001100110011001100,
64'b1100110011001100110011001100110000110011110011000011001111001100,
64'b0101010110101010010101011010101000000000000000000000000000000000,
64'b1001011010010110100101101001011010010110011010010110100110010110,
64'b1010010101011010101001010101101001101001100101100110100110010110,
64'b1100001100111100110000110011110001010101010101011010101010101010,
64'b1100001111000011001111000011110011110000000011110000111111110000,
64'b1010010110100101010110100101101010010110100101101001011010010110,
64'b1010010110100101010110100101101001011010010110100101101001011010,
64'b1010101010101010101010101010101011110000111100001111000011110000,
64'b0011001100110011110011001100110010101010101010101010101010101010,
64'b1010101001010101010101011010101001011010010110100101101001011010,
64'b0110100110010110011010011001011010101010101010101010101010101010,
64'b1111111100000000111111110000000011110000111100001111000011110000,
64'b0101101001011010010110100101101000001111000011111111000011110000,
64'b1010010110100101010110100101101000000000000000000000000000000000,
64'b1001100110011001011001100110011000111100110000111100001100111100,
64'b0011110011000011110000110011110010010110011010010110100110010110,
64'b0011110000111100001111000011110011001100110011001100110011001100,
64'b1010101010101010101010101010101010101010010101010101010110101010,
64'b0000000011111111111111110000000001101001100101100110100110010110,
64'b1001011010010110100101101001011000110011110011000011001111001100,
64'b0000111111110000000011111111000011111111000000001111111100000000,
64'b1111000011110000111100001111000001100110011001100110011001100110,
64'b1001100110011001011001100110011000110011110011000011001111001100,
64'b1001011001101001011010011001011011001100110011001100110011001100,
64'b1111111111111111000000000000000011111111000000001111111100000000,
64'b0011001111001100001100111100110011111111000000001111111100000000,
64'b0011001111001100001100111100110010101010101010101010101010101010,
64'b1001011010010110100101101001011011110000000011110000111111110000,
64'b0101101010100101101001010101101010010110011010010110100110010110,
64'b1010010101011010101001010101101001011010010110100101101001011010,
64'b1100110011001100110011001100110000110011001100111100110011001100,
64'b1111111111111111000000000000000010010110011010010110100110010110,
64'b0110100110010110011010011001011000001111000011111111000011110000,
64'b1111111100000000111111110000000000000000000000000000000000000000,
64'b0110011001100110011001100110011010010110100101101001011010010110,
64'b1100001100111100110000110011110000001111000011111111000011110000,
64'b0101101010100101101001010101101011110000111100001111000011110000,
64'b1010101001010101010101011010101011111111111111110000000000000000,
64'b0000111100001111111100001111000011111111111111110000000000000000,
64'b1001100110011001011001100110011011001100110011001100110011001100,
64'b1001100110011001011001100110011000000000111111111111111100000000,
64'b0011110011000011110000110011110010010110011010010110100110010110,
64'b1010101010101010101010101010101010011001011001101001100101100110,
64'b0101010110101010010101011010101011110000111100001111000011110000,
64'b1001100110011001011001100110011010010110011010010110100110010110,
64'b1001100110011001011001100110011001010101101010100101010110101010,
64'b0110100110010110011010011001011010101010101010101010101010101010,
64'b0000111111110000000011111111000011000011001111001100001100111100,
64'b0000111100001111111100001111000011111111000000001111111100000000,
64'b0000000011111111111111110000000001010101101010100101010110101010,
64'b1001100101100110100110010110011000000000000000000000000000000000,
64'b1111111100000000111111110000000010101010101010101010101010101010,
64'b0000000000000000000000000000000001011010010110100101101001011010,
64'b1100110000110011001100111100110011111111111111110000000000000000,
64'b1010101001010101010101011010101010010110011010010110100110010110,
64'b1010101001010101010101011010101001101001011010011001011010010110,
64'b1001011001101001011010011001011011111111000000001111111100000000,
64'b1010010110100101010110100101101000111100110000111100001100111100,
64'b1001100101100110100110010110011010011001100110010110011001100110,
64'b0000000000000000000000000000000011001100110011001100110011001100,
64'b1010101001010101010101011010101001101001011010011001011010010110,
64'b1111111100000000111111110000000000000000111111111111111100000000,
64'b0101010101010101101010101010101011111111111111110000000000000000,
64'b0110100101101001100101101001011000000000111111111111111100000000,
64'b1111111111111111000000000000000001100110011001100110011001100110,
64'b0000000000000000000000000000000010100101010110101010010101011010,
64'b0000111100001111111100001111000001011010101001011010010101011010,
64'b1001100110011001011001100110011001100110100110011001100101100110,
64'b1001100110011001011001100110011010100101101001010101101001011010,
64'b1001011001101001011010011001011011110000000011110000111111110000,
64'b1001100101100110100110010110011001101001100101100110100110010110,
64'b0110100101101001100101101001011010011001011001101001100101100110,
64'b0000000000000000000000000000000000110011110011000011001111001100,
64'b0000000011111111111111110000000001011010010110100101101001011010,
64'b1010101001010101010101011010101010101010010101010101010110101010,
64'b0000000000000000000000000000000001100110011001100110011001100110,
64'b0110100101101001100101101001011001010101101010100101010110101010,
64'b0000000000000000000000000000000000111100001111000011110000111100,
64'b0011110000111100001111000011110001011010101001011010010101011010,
64'b1010010110100101010110100101101010010110100101101001011010010110,
64'b0110011001100110011001100110011010011001100110010110011001100110,
64'b0101101010100101101001010101101001010101010101011010101010101010,
64'b0011001100110011110011001100110000001111000011111111000011110000,
64'b1111000011110000111100001111000000001111111100000000111111110000,
64'b1100110011001100110011001100110011001100001100110011001111001100,
64'b1100001100111100110000110011110010011001011001101001100101100110,
64'b0110011010011001100110010110011010011001011001101001100101100110,
64'b0110011010011001100110010110011000110011001100111100110011001100,
64'b0110011001100110011001100110011010010110100101101001011010010110,
64'b1100001111000011001111000011110000110011001100111100110011001100,
64'b0000000000000000000000000000000000001111111100000000111111110000,
64'b1001100101100110100110010110011011001100001100110011001111001100,
64'b0110100101101001100101101001011001101001100101100110100110010110,
64'b0110011001100110011001100110011000111100001111000011110000111100,
64'b0000000000000000000000000000000001100110011001100110011001100110,
64'b1111111100000000111111110000000001010101101010100101010110101010,
64'b1100110000110011001100111100110010101010010101010101010110101010,
64'b1111111100000000111111110000000000001111000011111111000011110000,
64'b0110011001100110011001100110011010010110100101101001011010010110,
64'b1100001111000011001111000011110001101001011010011001011010010110,
64'b0110100101101001100101101001011011110000111100001111000011110000,
64'b1001011010010110100101101001011001101001100101100110100110010110,
64'b0000111111110000000011111111000011110000111100001111000011110000,
64'b1010101010101010101010101010101010101010010101010101010110101010,
64'b1100001111000011001111000011110000001111000011111111000011110000,
64'b1100001100111100110000110011110010010110011010010110100110010110,
64'b1001011010010110100101101001011000001111111100000000111111110000,
64'b0000000000000000000000000000000000111100001111000011110000111100,
64'b1111111111111111000000000000000000110011001100111100110011001100,
64'b0000111100001111111100001111000000110011001100111100110011001100,
64'b0101010101010101101010101010101001010101101010100101010110101010,
64'b0011110000111100001111000011110001101001100101100110100110010110,
64'b1001011010010110100101101001011011110000111100001111000011110000,
64'b1001011010010110100101101001011010101010101010101010101010101010,
64'b1010010101011010101001010101101011110000000011110000111111110000,
64'b0000000000000000000000000000000011111111111111110000000000000000,
64'b0110011001100110011001100110011010011001100110010110011001100110,
64'b1001100101100110100110010110011011000011001111001100001100111100,
64'b0000000000000000000000000000000011001100110011001100110011001100,
64'b0011001111001100001100111100110001011010101001011010010101011010,
64'b1100110000110011001100111100110011000011110000110011110000111100,
64'b1010010101011010101001010101101001010101101010100101010110101010,
64'b1100110000110011001100111100110011000011110000110011110000111100,
64'b0110100110010110011010011001011010010110011010010110100110010110,
64'b1100110011001100110011001100110010101010101010101010101010101010,
64'b1111000011110000111100001111000011111111000000001111111100000000,
64'b0011110000111100001111000011110011001100110011001100110011001100,
64'b0000000011111111111111110000000000000000111111111111111100000000,
64'b0000000011111111111111110000000010101010101010101010101010101010,
64'b1001011010010110100101101001011010010110100101101001011010010110,
64'b0101010101010101101010101010101001011010101001011010010101011010,
64'b0101101010100101101001010101101011110000111100001111000011110000,
64'b1111111111111111000000000000000011001100001100110011001111001100,
64'b1100001100111100110000110011110010100101010110101010010101011010,
64'b1100001111000011001111000011110010011001100110010110011001100110,
64'b1001011010010110100101101001011000001111111100000000111111110000,
64'b1001100110011001011001100110011010010110011010010110100110010110,
64'b1001100101100110100110010110011001100110011001100110011001100110,
64'b1100110011001100110011001100110011111111111111110000000000000000,
64'b1111000011110000111100001111000011110000111100001111000011110000,
64'b0011001100110011110011001100110011111111111111110000000000000000,
64'b0101010110101010010101011010101001100110011001100110011001100110,
64'b1100001100111100110000110011110011000011001111001100001100111100,
64'b0101101001011010010110100101101011001100001100110011001111001100,
64'b0011110000111100001111000011110001010101101010100101010110101010,
64'b0101101001011010010110100101101000001111000011111111000011110000,
64'b1001011010010110100101101001011001100110100110011001100101100110,
64'b1010101010101010101010101010101000111100001111000011110000111100,
64'b1111000000001111000011111111000010101010010101010101010110101010,
64'b0011001111001100001100111100110000111100110000111100001100111100,
64'b1111111100000000111111110000000010010110100101101001011010010110,
64'b1111000011110000111100001111000010101010101010101010101010101010,
64'b1111111100000000111111110000000001010101101010100101010110101010,
64'b1111000011110000111100001111000000000000000000000000000000000000,
64'b1001100110011001011001100110011010010110100101101001011010010110,
64'b1111000000001111000011111111000011110000000011110000111111110000,
64'b0011001111001100001100111100110000001111000011111111000011110000,
64'b0000111111110000000011111111000010011001100110010110011001100110,
64'b0011001111001100001100111100110011111111000000001111111100000000,
64'b1100001100111100110000110011110001101001011010011001011010010110,
64'b1100110011001100110011001100110010100101010110101010010101011010,
64'b0000000011111111111111110000000000110011001100111100110011001100,
64'b1010010110100101010110100101101001011010101001011010010101011010,
64'b0000000000000000000000000000000001101001100101100110100110010110,
64'b1111111100000000111111110000000011001100110011001100110011001100,
64'b1111111111111111000000000000000000110011001100111100110011001100,
64'b1111111100000000111111110000000000000000000000000000000000000000,
64'b0011110000111100001111000011110011000011001111001100001100111100,
64'b1010101001010101010101011010101000000000111111111111111100000000,
64'b1010010110100101010110100101101001010101101010100101010110101010,
64'b0000000011111111111111110000000010010110100101101001011010010110,
64'b0000111100001111111100001111000001010101010101011010101010101010,
64'b1111000000001111000011111111000011000011001111001100001100111100,
64'b1111000011110000111100001111000001100110100110011001100101100110,
64'b1111111111111111000000000000000011110000111100001111000011110000,
64'b1001100101100110100110010110011001100110100110011001100101100110,
64'b1010101010101010101010101010101001101001100101100110100110010110,
64'b0101010101010101101010101010101001011010010110100101101001011010,
64'b0000000000000000000000000000000011110000111100001111000011110000,
64'b0101010101010101101010101010101010101010101010101010101010101010,
64'b0000111111110000000011111111000011110000000011110000111111110000,
64'b0011001100110011110011001100110011111111111111110000000000000000,
64'b1001100101100110100110010110011010011001100110010110011001100110,
64'b0101010101010101101010101010101011000011001111001100001100111100,
64'b0101010110101010010101011010101011001100110011001100110011001100,
64'b1010101001010101010101011010101001011010101001011010010101011010,
64'b0101010110101010010101011010101011000011110000110011110000111100,
64'b0000000000000000000000000000000001010101101010100101010110101010,
64'b0110100101101001100101101001011011000011110000110011110000111100,
64'b1100110011001100110011001100110001101001100101100110100110010110,
64'b1001011010010110100101101001011001101001100101100110100110010110,
64'b1111000011110000111100001111000011000011001111001100001100111100,
64'b1111000011110000111100001111000011110000111100001111000011110000,
64'b0101010101010101101010101010101010010110011010010110100110010110,
64'b1111111100000000111111110000000000111100110000111100001100111100,
64'b0000000000000000000000000000000001010101101010100101010110101010,
64'b0011001100110011110011001100110011110000000011110000111111110000,
64'b1010101001010101010101011010101011001100001100110011001111001100,
64'b1001100101100110100110010110011011110000111100001111000011110000,
64'b0011001111001100001100111100110010011001011001101001100101100110,
64'b0110100110010110011010011001011001011010101001011010010101011010,
64'b1111111100000000111111110000000010100101101001010101101001011010,
64'b1100001100111100110000110011110011000011001111001100001100111100,
64'b1111111100000000111111110000000010010110011010010110100110010110,
64'b0000111111110000000011111111000011110000000011110000111111110000,
64'b0000111111110000000011111111000011111111000000001111111100000000,
64'b1001100110011001011001100110011000111100110000111100001100111100,
64'b1010101001010101010101011010101001011010101001011010010101011010,
64'b0000000000000000000000000000000010011001100110010110011001100110,
64'b1100001111000011001111000011110000000000111111111111111100000000,
64'b0011001111001100001100111100110010100101101001010101101001011010,
64'b1111000000001111000011111111000001010101101010100101010110101010,
64'b0011110011000011110000110011110011000011110000110011110000111100,
64'b0101010101010101101010101010101011001100001100110011001111001100,
64'b0000000011111111111111110000000010011001011001101001100101100110,
64'b1100110011001100110011001100110010100101010110101010010101011010,
64'b0110100101101001100101101001011000111100110000111100001100111100,
64'b1111000000001111000011111111000010101010010101010101010110101010,
64'b1111000000001111000011111111000001010101010101011010101010101010,
64'b0110100101101001100101101001011011110000000011110000111111110000,
64'b0110011010011001100110010110011001100110100110011001100101100110,
64'b1010101010101010101010101010101010010110100101101001011010010110,
64'b0011110011000011110000110011110001010101010101011010101010101010,
64'b0000111111110000000011111111000010011001011001101001100101100110,
64'b1001100110011001011001100110011010011001100110010110011001100110,
64'b0110100101101001100101101001011000001111111100000000111111110000,
64'b0000111111110000000011111111000010100101101001010101101001011010,
64'b1010101001010101010101011010101001101001011010011001011010010110,
64'b1001100101100110100110010110011000110011110011000011001111001100,
64'b0110100110010110011010011001011001011010101001011010010101011010,
64'b1010101001010101010101011010101010011001100110010110011001100110,
64'b1010101001010101010101011010101001100110011001100110011001100110,
64'b0110100110010110011010011001011010101010010101010101010110101010,
64'b0110100101101001100101101001011001101001011010011001011010010110,
64'b0110011001100110011001100110011001101001100101100110100110010110,
64'b1111000000001111000011111111000011001100110011001100110011001100,
64'b1010101001010101010101011010101001101001011010011001011010010110,
64'b0011110000111100001111000011110000111100001111000011110000111100,
64'b0110100110010110011010011001011010101010010101010101010110101010,
64'b1010101001010101010101011010101000110011110011000011001111001100,
64'b0011001100110011110011001100110001101001100101100110100110010110,
64'b1001011010010110100101101001011001011010010110100101101001011010,
64'b0000000011111111111111110000000011001100001100110011001111001100,
64'b1100001111000011001111000011110010010110100101101001011010010110,
64'b0110100101101001100101101001011010010110100101101001011010010110,
64'b1100001100111100110000110011110000110011001100111100110011001100,
64'b0011110000111100001111000011110001101001100101100110100110010110,
64'b1001011010010110100101101001011010010110011010010110100110010110,
64'b0011001111001100001100111100110011110000111100001111000011110000,
64'b0011001111001100001100111100110011000011001111001100001100111100,
64'b0011110000111100001111000011110010100101010110101010010101011010,
64'b0000111100001111111100001111000000110011001100111100110011001100,
64'b0101101010100101101001010101101010100101101001010101101001011010,
64'b1010010101011010101001010101101000111100110000111100001100111100,
64'b1010101010101010101010101010101000110011110011000011001111001100,
64'b1100001111000011001111000011110000001111000011111111000011110000,
64'b0101010110101010010101011010101001101001100101100110100110010110,
64'b1001100101100110100110010110011011000011001111001100001100111100,
64'b0000111111110000000011111111000011110000111100001111000011110000,
64'b1111000011110000111100001111000010010110011010010110100110010110,
64'b1100001100111100110000110011110000111100110000111100001100111100,
64'b0011110000111100001111000011110001010101101010100101010110101010,
64'b1010010101011010101001010101101011110000000011110000111111110000,
64'b1001011010010110100101101001011011001100001100110011001111001100,
64'b1100110011001100110011001100110011110000111100001111000011110000,
64'b0000111100001111111100001111000010011001011001101001100101100110,
64'b1001100110011001011001100110011001011010101001011010010101011010,
64'b0000111111110000000011111111000001011010010110100101101001011010,
64'b0000111111110000000011111111000001101001100101100110100110010110,
64'b1001100110011001011001100110011001100110100110011001100101100110,
64'b1100001111000011001111000011110000000000111111111111111100000000,
64'b0000000011111111111111110000000010101010010101010101010110101010,
64'b1111111100000000111111110000000011000011110000110011110000111100,
64'b1111000000001111000011111111000001011010101001011010010101011010,
64'b0000111111110000000011111111000010101010101010101010101010101010,
64'b1100110000110011001100111100110010101010101010101010101010101010,
64'b1100001100111100110000110011110000111100110000111100001100111100,
64'b1111000011110000111100001111000001100110011001100110011001100110,
64'b1111111100000000111111110000000010101010010101010101010110101010,
64'b1001011010010110100101101001011000110011001100111100110011001100,
64'b0101010110101010010101011010101001011010010110100101101001011010,
64'b1001011001101001011010011001011000000000111111111111111100000000,
64'b1100110011001100110011001100110000110011001100111100110011001100,
64'b0101010110101010010101011010101010100101101001010101101001011010,
64'b0000000000000000000000000000000011001100110011001100110011001100,
64'b1010101001010101010101011010101001011010010110100101101001011010,
64'b0000000011111111111111110000000001100110100110011001100101100110,
64'b1001100101100110100110010110011001010101010101011010101010101010,
64'b1010010101011010101001010101101001100110100110011001100101100110,
64'b1100001111000011001111000011110001101001011010011001011010010110,
64'b1100110011001100110011001100110010100101010110101010010101011010,
64'b1001011001101001011010011001011001011010101001011010010101011010,
64'b0011110000111100001111000011110010100101010110101010010101011010,
64'b0000111111110000000011111111000001011010010110100101101001011010,
64'b0000000011111111111111110000000001010101010101011010101010101010,
64'b1010101010101010101010101010101001011010010110100101101001011010,
64'b1100001111000011001111000011110010011001011001101001100101100110,
64'b0101010101010101101010101010101001011010010110100101101001011010,
64'b1100110000110011001100111100110000110011110011000011001111001100,
64'b0101010101010101101010101010101011000011110000110011110000111100,
64'b0101101001011010010110100101101001100110011001100110011001100110,
64'b0110011001100110011001100110011001101001011010011001011010010110,
64'b1001011010010110100101101001011001101001100101100110100110010110,
64'b0110100110010110011010011001011001100110100110011001100101100110,
64'b0101010101010101101010101010101011001100001100110011001111001100,
64'b0101101001011010010110100101101001100110100110011001100101100110,
64'b0011110000111100001111000011110000110011110011000011001111001100,
64'b1111111111111111000000000000000011001100110011001100110011001100,
64'b0110011001100110011001100110011010011001011001101001100101100110,
64'b0000111111110000000011111111000011000011110000110011110000111100,
64'b0110011001100110011001100110011000110011110011000011001111001100,
64'b1010010110100101010110100101101000001111000011111111000011110000,
64'b0110011001100110011001100110011000001111111100000000111111110000,
64'b1001100101100110100110010110011010010110100101101001011010010110,
64'b0011110000111100001111000011110011000011001111001100001100111100,
64'b1100001100111100110000110011110010010110011010010110100110010110,
64'b0011110011000011110000110011110011000011110000110011110000111100,
64'b1100110011001100110011001100110010100101101001010101101001011010,
64'b1001100101100110100110010110011001101001011010011001011010010110,
64'b0000111111110000000011111111000001011010010110100101101001011010,
64'b1001011010010110100101101001011011001100110011001100110011001100,
64'b0110011001100110011001100110011000110011001100111100110011001100,
64'b1111000000001111000011111111000011111111000000001111111100000000,
64'b0110100101101001100101101001011011110000111100001111000011110000,
64'b1100110011001100110011001100110000000000000000000000000000000000,
64'b1001011010010110100101101001011010101010010101010101010110101010,
64'b1111000011110000111100001111000011110000000011110000111111110000,
64'b1010010110100101010110100101101001011010010110100101101001011010,
64'b0110100101101001100101101001011010100101101001010101101001011010,
64'b1100001111000011001111000011110010010110100101101001011010010110,
64'b0011001111001100001100111100110011110000111100001111000011110000,
64'b0011110011000011110000110011110010010110100101101001011010010110,
64'b0011110000111100001111000011110001011010010110100101101001011010,
64'b0101010110101010010101011010101011110000111100001111000011110000,
64'b1100110011001100110011001100110011110000111100001111000011110000,
64'b1111000000001111000011111111000001010101010101011010101010101010,
64'b0011110011000011110000110011110011111111000000001111111100000000,
64'b1010010101011010101001010101101000000000000000000000000000000000,
64'b1100001100111100110000110011110000110011001100111100110011001100,
64'b1100110000110011001100111100110010101010010101010101010110101010,
64'b1001100110011001011001100110011010011001011001101001100101100110,
64'b1111000011110000111100001111000000110011110011000011001111001100,
64'b1001011010010110100101101001011001101001100101100110100110010110,
64'b1100110000110011001100111100110011111111000000001111111100000000,
64'b0000111100001111111100001111000011000011001111001100001100111100,
64'b0110011001100110011001100110011000110011110011000011001111001100,
64'b0000111100001111111100001111000011111111000000001111111100000000,
64'b0000000000000000000000000000000011111111000000001111111100000000,
64'b1111000000001111000011111111000011001100110011001100110011001100,
64'b0000111111110000000011111111000001010101010101011010101010101010,
64'b1001100110011001011001100110011000000000000000000000000000000000,
64'b1111000000001111000011111111000011110000111100001111000011110000,
64'b0011110000111100001111000011110010011001100110010110011001100110,
64'b0011110011000011110000110011110001101001011010011001011010010110,
64'b1100110011001100110011001100110000001111000011111111000011110000,
64'b1111000011110000111100001111000000111100110000111100001100111100,
64'b0110011010011001100110010110011011111111111111110000000000000000,
64'b1010101010101010101010101010101011110000000011110000111111110000,
64'b0101010110101010010101011010101011110000111100001111000011110000,
64'b0101010110101010010101011010101011111111111111110000000000000000,
64'b1010101010101010101010101010101011111111111111110000000000000000,
64'b0000000011111111111111110000000011110000111100001111000011110000,
64'b1010101001010101010101011010101011001100110011001100110011001100,
64'b0011110000111100001111000011110010101010101010101010101010101010,
64'b1010101001010101010101011010101011111111000000001111111100000000,
64'b1010010101011010101001010101101000111100001111000011110000111100,
64'b1111000000001111000011111111000001101001100101100110100110010110,
64'b0101101001011010010110100101101001010101101010100101010110101010,
64'b1111111100000000111111110000000001011010101001011010010101011010,
64'b1100001111000011001111000011110010101010101010101010101010101010,
64'b0110011001100110011001100110011010101010010101010101010110101010,
64'b1100110011001100110011001100110001010101101010100101010110101010,
64'b0011001100110011110011001100110010101010101010101010101010101010,
64'b1100110011001100110011001100110010101010101010101010101010101010,
64'b1111111111111111000000000000000001010101101010100101010110101010,
64'b1001100110011001011001100110011011110000111100001111000011110000,
64'b1010010101011010101001010101101011001100110011001100110011001100,
64'b0011001100110011110011001100110011111111111111110000000000000000,
64'b0110011010011001100110010110011000001111111100000000111111110000,
64'b0000000011111111111111110000000000111100110000111100001100111100,
64'b1001100101100110100110010110011000110011001100111100110011001100,
64'b1111111111111111000000000000000011001100001100110011001111001100,
64'b0000111111110000000011111111000001100110011001100110011001100110,
64'b1001011010010110100101101001011000110011001100111100110011001100,
64'b1111000011110000111100001111000001100110011001100110011001100110,
64'b1111000011110000111100001111000001100110011001100110011001100110,
64'b0101101001011010010110100101101011001100110011001100110011001100,
64'b0000000000000000000000000000000000110011001100111100110011001100,
64'b1001011010010110100101101001011011111111000000001111111100000000,
64'b0110011010011001100110010110011011110000111100001111000011110000,
64'b1111000011110000111100001111000000000000000000000000000000000000,
64'b0110100101101001100101101001011010101010010101010101010110101010,
64'b0101010101010101101010101010101011110000000011110000111111110000,
64'b0110100101101001100101101001011001011010010110100101101001011010,
64'b0000000000000000000000000000000010100101101001010101101001011010,
64'b1010101001010101010101011010101010010110100101101001011010010110,
64'b1100001100111100110000110011110011110000111100001111000011110000,
64'b1111111100000000111111110000000010010110100101101001011010010110,
64'b0000111100001111111100001111000001011010101001011010010101011010,
64'b0000111111110000000011111111000000000000000000000000000000000000,
64'b0101101010100101101001010101101000000000000000000000000000000000,
64'b0110011010011001100110010110011001100110011001100110011001100110,
64'b1010010110100101010110100101101001010101101010100101010110101010,
64'b1010010101011010101001010101101001100110100110011001100101100110,
64'b0011001100110011110011001100110000000000111111111111111100000000,
64'b0101101010100101101001010101101011000011001111001100001100111100,
64'b0011110000111100001111000011110000111100001111000011110000111100,
64'b0110100110010110011010011001011000001111111100000000111111110000,
64'b1100001111000011001111000011110000001111000011111111000011110000,
64'b1111111100000000111111110000000001101001011010011001011010010110,
64'b1111000011110000111100001111000011110000111100001111000011110000,
64'b0101101010100101101001010101101001100110100110011001100101100110,
64'b1010010110100101010110100101101010101010101010101010101010101010,
64'b1001011010010110100101101001011000000000000000000000000000000000,
64'b0000111111110000000011111111000000111100001111000011110000111100,
64'b0011110011000011110000110011110000110011001100111100110011001100,
64'b1100001111000011001111000011110011000011110000110011110000111100,
64'b1100001111000011001111000011110001010101010101011010101010101010,
64'b0011110000111100001111000011110001011010101001011010010101011010,
64'b1001100101100110100110010110011000001111111100000000111111110000,
64'b0101010101010101101010101010101000000000111111111111111100000000,
64'b1100110000110011001100111100110011111111000000001111111100000000,
64'b1010101001010101010101011010101001101001100101100110100110010110,
64'b0000111111110000000011111111000001010101101010100101010110101010,
64'b1100001100111100110000110011110001101001011010011001011010010110,
64'b1001011010010110100101101001011001100110011001100110011001100110,
64'b0011001100110011110011001100110000000000000000000000000000000000,
64'b0110011001100110011001100110011000001111111100000000111111110000,
64'b0101010110101010010101011010101011110000111100001111000011110000,
64'b0000000000000000000000000000000010100101010110101010010101011010,
64'b1001011001101001011010011001011001100110011001100110011001100110,
64'b1111111111111111000000000000000001100110100110011001100101100110,
64'b1111111111111111000000000000000010101010010101010101010110101010,
64'b1010010101011010101001010101101011111111111111110000000000000000,
64'b0110011001100110011001100110011001010101010101011010101010101010,
64'b0110011010011001100110010110011000111100110000111100001100111100,
64'b1010010101011010101001010101101011001100110011001100110011001100,
64'b0101101010100101101001010101101001101001100101100110100110010110,
64'b1100001100111100110000110011110010010110100101101001011010010110,
64'b1111000011110000111100001111000000000000000000000000000000000000,
64'b1001011010010110100101101001011000000000111111111111111100000000,
64'b0011001100110011110011001100110011111111000000001111111100000000,
64'b0000000000000000000000000000000011001100001100110011001111001100,
64'b0011110011000011110000110011110000111100001111000011110000111100,
64'b1010101010101010101010101010101011000011110000110011110000111100,
64'b1010101010101010101010101010101010011001100110010110011001100110,
64'b0110011010011001100110010110011010101010101010101010101010101010,
64'b0011110000111100001111000011110001100110011001100110011001100110,
64'b1100001111000011001111000011110001011010101001011010010101011010,
64'b1001100101100110100110010110011001011010010110100101101001011010,
64'b1100001100111100110000110011110000111100110000111100001100111100,
64'b0101010101010101101010101010101011000011001111001100001100111100,
64'b1010010110100101010110100101101000000000000000000000000000000000,
64'b1010010110100101010110100101101011111111111111110000000000000000,
64'b0101010101010101101010101010101001010101010101011010101010101010,
64'b0000111111110000000011111111000000001111000011111111000011110000,
64'b1100001100111100110000110011110010100101010110101010010101011010,
64'b0011110011000011110000110011110000001111111100000000111111110000,
64'b1111000011110000111100001111000010010110100101101001011010010110,
64'b1010101001010101010101011010101001100110011001100110011001100110,
64'b0110011010011001100110010110011000111100001111000011110000111100,
64'b1111000011110000111100001111000011001100001100110011001111001100,
64'b0110011001100110011001100110011010011001011001101001100101100110,
64'b1111111100000000111111110000000001011010101001011010010101011010,
64'b1100001100111100110000110011110001011010101001011010010101011010,
64'b1100001111000011001111000011110000000000000000000000000000000000,
64'b1111111111111111000000000000000000000000000000000000000000000000,
64'b1100001111000011001111000011110001100110011001100110011001100110,
64'b0000111100001111111100001111000001010101101010100101010110101010,
64'b1100001100111100110000110011110001100110100110011001100101100110,
64'b1010101010101010101010101010101000000000111111111111111100000000,
64'b0110100110010110011010011001011011000011001111001100001100111100,
64'b0101101010100101101001010101101000111100001111000011110000111100,
64'b1010101010101010101010101010101000001111111100000000111111110000,
64'b1010101010101010101010101010101000001111000011111111000011110000,
64'b1100110011001100110011001100110010010110100101101001011010010110,
64'b0101010101010101101010101010101011000011001111001100001100111100,
64'b1111000000001111000011111111000001101001011010011001011010010110,
64'b0000111111110000000011111111000011110000000011110000111111110000,
64'b1010101010101010101010101010101001100110100110011001100101100110,
64'b1010010101011010101001010101101010011001100110010110011001100110,
64'b0101010110101010010101011010101010010110011010010110100110010110,
64'b0101101010100101101001010101101011110000111100001111000011110000,
64'b1100110011001100110011001100110000001111111100000000111111110000,
64'b0011110011000011110000110011110001100110100110011001100101100110,
64'b1100110000110011001100111100110001100110011001100110011001100110,
64'b0110011001100110011001100110011011000011001111001100001100111100,
64'b1100110011001100110011001100110000000000000000000000000000000000,
64'b1111000011110000111100001111000010011001011001101001100101100110,
64'b0110100101101001100101101001011011111111000000001111111100000000,
64'b1010010110100101010110100101101011001100110011001100110011001100,
64'b1111000011110000111100001111000011110000111100001111000011110000,
64'b1010101001010101010101011010101000001111111100000000111111110000,
64'b0110100110010110011010011001011000110011001100111100110011001100,
64'b1001011001101001011010011001011000110011001100111100110011001100,
64'b1111111100000000111111110000000001100110100110011001100101100110,
64'b0000000011111111111111110000000001011010010110100101101001011010,
64'b1100110000110011001100111100110011111111111111110000000000000000,
64'b1100110000110011001100111100110011111111000000001111111100000000,
64'b0101010101010101101010101010101000110011110011000011001111001100,
64'b0000111111110000000011111111000011111111000000001111111100000000,
64'b0000111111110000000011111111000011001100110011001100110011001100,
64'b0110011010011001100110010110011011111111111111110000000000000000,
64'b1001011010010110100101101001011011110000111100001111000011110000,
64'b0000111100001111111100001111000011111111000000001111111100000000,
64'b0101010110101010010101011010101000000000111111111111111100000000,
64'b0011001111001100001100111100110011110000111100001111000011110000,
64'b1001100110011001011001100110011001011010010110100101101001011010,
64'b0110011001100110011001100110011001101001011010011001011010010110,
64'b1010010101011010101001010101101010011001011001101001100101100110,
64'b1001100110011001011001100110011000000000000000000000000000000000,
64'b1100110000110011001100111100110001010101010101011010101010101010,
64'b1010010110100101010110100101101000001111000011111111000011110000,
64'b0101010101010101101010101010101011111111111111110000000000000000,
64'b0000111111110000000011111111000011110000111100001111000011110000,
64'b1100001111000011001111000011110010101010101010101010101010101010,
64'b0110100110010110011010011001011001010101101010100101010110101010,
64'b1111111100000000111111110000000011111111111111110000000000000000,
64'b1001100110011001011001100110011011111111111111110000000000000000,
64'b0000111100001111111100001111000001010101101010100101010110101010,
64'b0011110000111100001111000011110000110011110011000011001111001100,
64'b1001011010010110100101101001011011000011001111001100001100111100,
64'b1100110000110011001100111100110001101001011010011001011010010110,
64'b0011110000111100001111000011110000000000000000000000000000000000,
64'b1010010110100101010110100101101011001100110011001100110011001100,
64'b1001100101100110100110010110011001010101101010100101010110101010,
64'b0110011001100110011001100110011010101010101010101010101010101010,
64'b0101010110101010010101011010101001010101101010100101010110101010,
64'b1010101001010101010101011010101011000011110000110011110000111100,
64'b1001100110011001011001100110011000111100110000111100001100111100,
64'b1010010101011010101001010101101001011010101001011010010101011010,
64'b0101101010100101101001010101101011001100001100110011001111001100,
64'b1111000000001111000011111111000000111100001111000011110000111100,
64'b0000000000000000000000000000000010101010010101010101010110101010,
64'b1111000000001111000011111111000011000011001111001100001100111100,
64'b0101010110101010010101011010101010011001100110010110011001100110,
64'b1001100101100110100110010110011010010110100101101001011010010110,
64'b0101101001011010010110100101101010011001011001101001100101100110,
64'b1010101010101010101010101010101011110000111100001111000011110000,
64'b1100001100111100110000110011110000110011110011000011001111001100,
64'b0011110000111100001111000011110000111100001111000011110000111100,
64'b0011110000111100001111000011110000001111111100000000111111110000,
64'b1001100101100110100110010110011001011010101001011010010101011010,
64'b0011110000111100001111000011110001100110100110011001100101100110,
64'b1010101010101010101010101010101010100101101001010101101001011010,
64'b0000111111110000000011111111000010100101010110101010010101011010,
64'b0000111111110000000011111111000000110011001100111100110011001100,
64'b0011001111001100001100111100110001011010101001011010010101011010,
64'b1100001100111100110000110011110000111100001111000011110000111100,
64'b1111111111111111000000000000000001101001100101100110100110010110,
64'b0101101001011010010110100101101011000011110000110011110000111100,
64'b0000111100001111111100001111000011111111000000001111111100000000,
64'b0000111100001111111100001111000000001111000011111111000011110000,
64'b1111111100000000111111110000000000001111111100000000111111110000,
64'b0000000011111111111111110000000010101010010101010101010110101010,
64'b1100110000110011001100111100110011001100001100110011001111001100,
64'b0101010101010101101010101010101001101001011010011001011010010110,
64'b1010101001010101010101011010101010011001011001101001100101100110,
64'b1010010101011010101001010101101001100110100110011001100101100110,
64'b1010010110100101010110100101101011110000111100001111000011110000,
64'b0011110000111100001111000011110001100110100110011001100101100110,
64'b1010101010101010101010101010101010100101010110101010010101011010,
64'b0011110000111100001111000011110000111100110000111100001100111100,
64'b1111000011110000111100001111000000001111111100000000111111110000,
64'b0011110011000011110000110011110001010101010101011010101010101010,
64'b1010101010101010101010101010101011111111000000001111111100000000,
64'b0101101001011010010110100101101001010101101010100101010110101010,
64'b0101010101010101101010101010101000110011001100111100110011001100,
64'b1010010110100101010110100101101010100101101001010101101001011010,
64'b0110011001100110011001100110011001101001100101100110100110010110,
64'b1001100110011001011001100110011001101001011010011001011010010110,
64'b0110011010011001100110010110011011000011110000110011110000111100,
64'b0011001111001100001100111100110001010101101010100101010110101010,
64'b1010010101011010101001010101101011000011110000110011110000111100,
64'b1100110011001100110011001100110001100110100110011001100101100110,
64'b0000111111110000000011111111000011110000000011110000111111110000,
64'b1111111100000000111111110000000010101010010101010101010110101010,
64'b1111000000001111000011111111000011001100110011001100110011001100,
64'b0110011001100110011001100110011001010101010101011010101010101010,
64'b0011001111001100001100111100110011001100110011001100110011001100,
64'b1100110011001100110011001100110001011010010110100101101001011010,
64'b1001100101100110100110010110011010011001011001101001100101100110,
64'b1001011010010110100101101001011010010110011010010110100110010110,
64'b0011110000111100001111000011110011000011001111001100001100111100,
64'b0110100101101001100101101001011010100101010110101010010101011010,
64'b1010010110100101010110100101101010011001100110010110011001100110,
64'b1100110000110011001100111100110000001111111100000000111111110000,
64'b1111000011110000111100001111000001101001011010011001011010010110,
64'b0000000011111111111111110000000010101010010101010101010110101010,
64'b1111111111111111000000000000000010011001100110010110011001100110,
64'b0000000011111111111111110000000001011010010110100101101001011010,
64'b1001011010010110100101101001011011001100110011001100110011001100,
64'b1111000011110000111100001111000001011010010110100101101001011010,
64'b1111000011110000111100001111000000110011110011000011001111001100,
64'b1100001111000011001111000011110011000011110000110011110000111100,
64'b1100001100111100110000110011110000111100110000111100001100111100,
64'b0000111111110000000011111111000001011010101001011010010101011010,
64'b1100001100111100110000110011110011001100001100110011001111001100,
64'b1001100101100110100110010110011000111100001111000011110000111100,
64'b1010010110100101010110100101101010101010010101010101010110101010,
64'b0101010110101010010101011010101011000011001111001100001100111100,
64'b1111111111111111000000000000000010011001100110010110011001100110,
64'b1010101010101010101010101010101010010110100101101001011010010110,
64'b0101010101010101101010101010101010011001011001101001100101100110,
64'b0110100110010110011010011001011011110000111100001111000011110000,
64'b1111111100000000111111110000000000110011110011000011001111001100,
64'b1010101001010101010101011010101011110000000011110000111111110000,
64'b1111111111111111000000000000000010101010101010101010101010101010,
64'b0011110000111100001111000011110001101001100101100110100110010110,
64'b1010010101011010101001010101101000001111111100000000111111110000,
64'b0000111111110000000011111111000001010101101010100101010110101010,
64'b1010010101011010101001010101101011110000000011110000111111110000,
64'b0000000011111111111111110000000000001111111100000000111111110000,
64'b0101010110101010010101011010101010100101101001010101101001011010,
64'b0110100110010110011010011001011010011001100110010110011001100110,
64'b1100110000110011001100111100110011001100110011001100110011001100,
64'b1100001111000011001111000011110000001111111100000000111111110000,
64'b0101101010100101101001010101101010100101010110101010010101011010,
64'b0110011001100110011001100110011011111111000000001111111100000000,
64'b1001100101100110100110010110011000000000111111111111111100000000,
64'b0101010101010101101010101010101001100110011001100110011001100110,
64'b1001100101100110100110010110011000111100110000111100001100111100,
64'b0110100101101001100101101001011000000000111111111111111100000000,
64'b0000111100001111111100001111000000110011001100111100110011001100,
64'b0110100101101001100101101001011000000000111111111111111100000000,
64'b1111111100000000111111110000000010101010010101010101010110101010,
64'b1100110000110011001100111100110000110011110011000011001111001100,
64'b0101010101010101101010101010101010010110100101101001011010010110,
64'b1100001100111100110000110011110001011010010110100101101001011010,
64'b0110011010011001100110010110011000000000111111111111111100000000,
64'b0011110000111100001111000011110011001100001100110011001111001100,
64'b1111000011110000111100001111000000000000000000000000000000000000,
64'b1100001100111100110000110011110001010101010101011010101010101010,
64'b0011001100110011110011001100110010010110100101101001011010010110,
64'b0101010101010101101010101010101011110000000011110000111111110000,
64'b0110011001100110011001100110011001010101010101011010101010101010,
64'b0101101001011010010110100101101001011010010110100101101001011010,
64'b1100110011001100110011001100110001010101010101011010101010101010,
64'b0101010110101010010101011010101010011001100110010110011001100110,
64'b0101101010100101101001010101101010100101101001010101101001011010,
64'b0000111111110000000011111111000011000011001111001100001100111100,
64'b1001011010010110100101101001011000110011110011000011001111001100,
64'b0000000000000000000000000000000011111111111111110000000000000000,
64'b1111111111111111000000000000000010100101101001010101101001011010,
64'b1001100101100110100110010110011010101010101010101010101010101010,
64'b0101101010100101101001010101101011001100110011001100110011001100,
64'b1111000011110000111100001111000001101001100101100110100110010110,
64'b0110011001100110011001100110011000000000111111111111111100000000,
64'b1001011010010110100101101001011001100110011001100110011001100110,
64'b0011001111001100001100111100110010011001011001101001100101100110,
64'b1111000011110000111100001111000011001100110011001100110011001100,
64'b0011001100110011110011001100110010010110100101101001011010010110,
64'b1100110000110011001100111100110010011001011001101001100101100110,
64'b1010101001010101010101011010101001011010101001011010010101011010,
64'b1100001100111100110000110011110000001111000011111111000011110000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000010011001011001101001100101100110,
64'b1001011010010110100101101001011001100110011001100110011001100110,
64'b1100110011001100110011001100110011110000111100001111000011110000,
64'b1010101001010101010101011010101000111100110000111100001100111100,
64'b0000000000000000000000000000000011111111111111110000000000000000,
64'b0110011001100110011001100110011010010110100101101001011010010110,
64'b0000000011111111111111110000000011000011110000110011110000111100,
64'b0101101001011010010110100101101011110000111100001111000011110000,
64'b1111000000001111000011111111000011000011001111001100001100111100,
64'b1111000000001111000011111111000011000011110000110011110000111100,
64'b1111000000001111000011111111000011001100001100110011001111001100,
64'b1001011010010110100101101001011001010101101010100101010110101010,
64'b1100001111000011001111000011110010101010101010101010101010101010,
64'b0101101010100101101001010101101011000011110000110011110000111100,
64'b1010010101011010101001010101101000111100001111000011110000111100,
64'b0101101010100101101001010101101001010101101010100101010110101010,
64'b1100110011001100110011001100110011110000000011110000111111110000,
64'b1001011010010110100101101001011010101010101010101010101010101010,
64'b1001100101100110100110010110011001101001100101100110100110010110,
64'b1111000000001111000011111111000000001111111100000000111111110000,
64'b0011110000111100001111000011110001010101101010100101010110101010,
64'b0000000000000000000000000000000011110000000011110000111111110000,
64'b1111111111111111000000000000000000001111111100000000111111110000,
64'b1100001111000011001111000011110010100101101001010101101001011010,
64'b1010010110100101010110100101101010011001100110010110011001100110,
64'b1100110000110011001100111100110011001100110011001100110011001100,
64'b0011110000111100001111000011110000001111111100000000111111110000,
64'b1111111100000000111111110000000010100101010110101010010101011010,
64'b1100110000110011001100111100110010011001011001101001100101100110,
64'b0101101001011010010110100101101011111111000000001111111100000000,
64'b1100001100111100110000110011110001011010010110100101101001011010,
64'b1100001111000011001111000011110010011001100110010110011001100110,
64'b0000000011111111111111110000000000001111000011111111000011110000,
64'b1010010101011010101001010101101010010110011010010110100110010110,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000011111111111111110000000000000000,
64'b1010010101011010101001010101101001011010010110100101101001011010,
64'b1001100101100110100110010110011001011010101001011010010101011010,
64'b1010010110100101010110100101101010011001100110010110011001100110,
64'b1010010101011010101001010101101001011010010110100101101001011010,
64'b0000000000000000000000000000000001010101101010100101010110101010,
64'b1010010101011010101001010101101011000011001111001100001100111100,
64'b0110011010011001100110010110011000000000000000000000000000000000,
64'b1100110000110011001100111100110000001111111100000000111111110000,
64'b1010101010101010101010101010101010011001011001101001100101100110,
64'b0101101010100101101001010101101001011010010110100101101001011010,
64'b1100001111000011001111000011110000110011001100111100110011001100,
64'b0000000011111111111111110000000010101010010101010101010110101010,
64'b0101010110101010010101011010101001010101101010100101010110101010,
64'b1010010110100101010110100101101011110000111100001111000011110000,
64'b0000111111110000000011111111000000000000000000000000000000000000,
64'b1111000000001111000011111111000001010101010101011010101010101010,
64'b0011110000111100001111000011110011000011110000110011110000111100,
64'b0110011001100110011001100110011010101010101010101010101010101010,
64'b1100110011001100110011001100110011110000000011110000111111110000,
64'b0011110000111100001111000011110000000000000000000000000000000000,
64'b1001100110011001011001100110011000000000111111111111111100000000,
64'b1100001100111100110000110011110011000011110000110011110000111100,
64'b1100001111000011001111000011110000110011110011000011001111001100,
64'b0000000000000000000000000000000011110000111100001111000011110000,
64'b0101010110101010010101011010101010011001100110010110011001100110,
64'b1100110000110011001100111100110010011001100110010110011001100110,
64'b0101101001011010010110100101101011111111000000001111111100000000,
64'b0110011001100110011001100110011000000000000000000000000000000000,
64'b1100001100111100110000110011110011001100110011001100110011001100,
64'b1111111111111111000000000000000010100101010110101010010101011010,
64'b0101101001011010010110100101101001100110011001100110011001100110,
64'b0101101001011010010110100101101000000000111111111111111100000000,
64'b0000111111110000000011111111000010101010101010101010101010101010,
64'b0011110000111100001111000011110011111111111111110000000000000000,
64'b0101101010100101101001010101101010100101010110101010010101011010,
64'b0000111111110000000011111111000010100101101001010101101001011010,
64'b1010101010101010101010101010101011111111000000001111111100000000,
64'b0011001100110011110011001100110000111100001111000011110000111100,
64'b0000111100001111111100001111000010010110100101101001011010010110,
64'b1001100101100110100110010110011001010101010101011010101010101010,
64'b0011110000111100001111000011110000000000000000000000000000000000,
64'b1111000000001111000011111111000011110000111100001111000011110000,
64'b0000000000000000000000000000000011001100001100110011001111001100,
64'b1001100101100110100110010110011000111100001111000011110000111100,
64'b0011001100110011110011001100110011111111000000001111111100000000,
64'b1111111100000000111111110000000010011001100110010110011001100110,
64'b0011001111001100001100111100110000111100001111000011110000111100,
64'b0110100101101001100101101001011011000011110000110011110000111100,
64'b1010010110100101010110100101101000111100001111000011110000111100,
64'b0110100110010110011010011001011011110000000011110000111111110000,
64'b1111000000001111000011111111000000001111000011111111000011110000,
64'b0000000000000000000000000000000010010110100101101001011010010110,
64'b0000000011111111111111110000000010100101010110101010010101011010,
64'b1100001111000011001111000011110001100110100110011001100101100110,
64'b1100001100111100110000110011110000111100110000111100001100111100,
64'b1111000000001111000011111111000001010101101010100101010110101010,
64'b0101101001011010010110100101101011000011001111001100001100111100,
64'b0101101010100101101001010101101011111111111111110000000000000000,
64'b1010101010101010101010101010101000111100001111000011110000111100,
64'b0011001100110011110011001100110010100101010110101010010101011010,
64'b0110011001100110011001100110011000001111111100000000111111110000,
64'b1001011010010110100101101001011010100101010110101010010101011010,
64'b0011001100110011110011001100110000000000111111111111111100000000,
64'b0000000000000000000000000000000001010101101010100101010110101010,
64'b1111111100000000111111110000000001101001100101100110100110010110,
64'b1001011001101001011010011001011011001100001100110011001111001100,
64'b0110100101101001100101101001011011000011110000110011110000111100,
64'b1001100101100110100110010110011001011010101001011010010101011010,
64'b0101101001011010010110100101101010011001100110010110011001100110,
64'b1111111100000000111111110000000000001111111100000000111111110000,
64'b1100110011001100110011001100110010101010101010101010101010101010,
64'b1001100110011001011001100110011010100101010110101010010101011010,
64'b1100110011001100110011001100110011001100001100110011001111001100,
64'b0011001111001100001100111100110000000000111111111111111100000000,
64'b1100110011001100110011001100110011001100001100110011001111001100,
64'b0101010110101010010101011010101011111111111111110000000000000000,
64'b1010101001010101010101011010101010011001100110010110011001100110,
64'b1010101001010101010101011010101000111100110000111100001100111100,
64'b0101010101010101101010101010101000001111000011111111000011110000,
64'b1010010110100101010110100101101010100101010110101010010101011010,
64'b1010101010101010101010101010101001100110100110011001100101100110,
64'b0110100101101001100101101001011010010110100101101001011010010110,
64'b0110011001100110011001100110011001010101101010100101010110101010,
64'b1111000011110000111100001111000001100110011001100110011001100110,
64'b0011110000111100001111000011110011001100001100110011001111001100,
64'b0101101001011010010110100101101000001111000011111111000011110000,
64'b0000111100001111111100001111000001010101010101011010101010101010,
64'b1111000011110000111100001111000010100101101001010101101001011010,
64'b0011001100110011110011001100110010101010101010101010101010101010,
64'b0011001100110011110011001100110010010110100101101001011010010110,
64'b1001100110011001011001100110011001011010101001011010010101011010,
64'b0110011001100110011001100110011001010101101010100101010110101010,
64'b1001100101100110100110010110011001100110100110011001100101100110,
64'b0110011001100110011001100110011011000011110000110011110000111100,
64'b1100001100111100110000110011110001101001100101100110100110010110,
64'b1001011010010110100101101001011011001100110011001100110011001100,
64'b0101010110101010010101011010101000111100001111000011110000111100,
64'b0000111111110000000011111111000000001111000011111111000011110000,
64'b0011001111001100001100111100110001010101101010100101010110101010,
64'b1111111100000000111111110000000001100110011001100110011001100110,
64'b0101010110101010010101011010101010011001011001101001100101100110,
64'b1111000011110000111100001111000001100110011001100110011001100110,
64'b0101101001011010010110100101101011000011001111001100001100111100,
64'b1001011010010110100101101001011011001100001100110011001111001100,
64'b1001011010010110100101101001011010011001100110010110011001100110,
64'b1100001111000011001111000011110011000011110000110011110000111100,
64'b0011110000111100001111000011110010100101010110101010010101011010,
64'b1111000000001111000011111111000010010110011010010110100110010110,
64'b1100001100111100110000110011110011110000111100001111000011110000,
64'b0011001100110011110011001100110000001111111100000000111111110000,
64'b0000000011111111111111110000000011111111000000001111111100000000,
64'b0000111100001111111100001111000010011001100110010110011001100110,
64'b1111111111111111000000000000000000111100001111000011110000111100,
64'b0011001100110011110011001100110011000011110000110011110000111100,
64'b1111111100000000111111110000000000111100001111000011110000111100,
64'b0011001111001100001100111100110011110000000011110000111111110000,
64'b1100001100111100110000110011110000001111000011111111000011110000,
64'b1100001100111100110000110011110010010110100101101001011010010110,
64'b0000111111110000000011111111000010100101010110101010010101011010,
64'b1010010101011010101001010101101001100110100110011001100101100110,
64'b0000000011111111111111110000000000111100110000111100001100111100,
64'b1010010101011010101001010101101001010101101010100101010110101010,
64'b1010101001010101010101011010101011001100001100110011001111001100,
64'b1001100110011001011001100110011000111100110000111100001100111100,
64'b0110011001100110011001100110011010101010101010101010101010101010,
64'b0000000011111111111111110000000010010110100101101001011010010110,
64'b0110100110010110011010011001011000111100110000111100001100111100,
64'b0000000011111111111111110000000000000000111111111111111100000000,
64'b1100001111000011001111000011110011001100110011001100110011001100,
64'b0101101001011010010110100101101010101010010101010101010110101010,
64'b0110100101101001100101101001011001101001100101100110100110010110,
64'b1111000000001111000011111111000000000000111111111111111100000000,
64'b0110100101101001100101101001011000001111111100000000111111110000,
64'b0011001100110011110011001100110010101010010101010101010110101010,
64'b0101010110101010010101011010101011001100110011001100110011001100,
64'b1001100101100110100110010110011010100101101001010101101001011010,
64'b0000111100001111111100001111000001011010101001011010010101011010,
64'b1111000011110000111100001111000001100110011001100110011001100110,
64'b1111111100000000111111110000000011000011001111001100001100111100,
64'b1111111111111111000000000000000011110000000011110000111111110000,
64'b1111111100000000111111110000000001010101010101011010101010101010,
64'b0110011010011001100110010110011001011010010110100101101001011010,
64'b1100001100111100110000110011110000110011001100111100110011001100,
64'b1010101001010101010101011010101010010110011010010110100110010110,
64'b0101101001011010010110100101101011111111111111110000000000000000,
64'b0000000011111111111111110000000010101010010101010101010110101010,
64'b0110100101101001100101101001011000110011001100111100110011001100,
64'b0011001111001100001100111100110001011010010110100101101001011010,
64'b0110100110010110011010011001011000110011110011000011001111001100,
64'b0110011010011001100110010110011001100110100110011001100101100110,
64'b0011001111001100001100111100110010010110100101101001011010010110,
64'b1111111100000000111111110000000011110000000011110000111111110000,
64'b0110100110010110011010011001011000000000111111111111111100000000,
64'b0101010110101010010101011010101001100110011001100110011001100110,
64'b0000000000000000000000000000000010011001011001101001100101100110,
64'b0000000011111111111111110000000011110000111100001111000011110000,
64'b0101101001011010010110100101101010010110011010010110100110010110,
64'b0110100101101001100101101001011010101010101010101010101010101010,
64'b1001011010010110100101101001011010011001100110010110011001100110,
64'b0101101010100101101001010101101001011010010110100101101001011010,
64'b0000111111110000000011111111000010011001011001101001100101100110,
64'b1001011001101001011010011001011000001111000011111111000011110000,
64'b1100001111000011001111000011110011000011110000110011110000111100,
64'b1010010110100101010110100101101001101001100101100110100110010110,
64'b1111111111111111000000000000000000000000111111111111111100000000,
64'b0011110011000011110000110011110001010101010101011010101010101010,
64'b0011001100110011110011001100110010010110100101101001011010010110,
64'b0000000000000000000000000000000011000011110000110011110000111100,
64'b1111111111111111000000000000000011111111000000001111111100000000,
64'b1001100101100110100110010110011000111100110000111100001100111100,
64'b1100001100111100110000110011110001100110011001100110011001100110,
64'b0110100110010110011010011001011000111100001111000011110000111100,
64'b1100110000110011001100111100110010011001011001101001100101100110,
64'b0101010110101010010101011010101000111100001111000011110000111100,
64'b1001011010010110100101101001011011111111000000001111111100000000,
64'b0011110011000011110000110011110010100101010110101010010101011010,
64'b1111111100000000111111110000000010010110011010010110100110010110,
64'b1010101001010101010101011010101011111111111111110000000000000000,
64'b0011001100110011110011001100110001100110011001100110011001100110,
64'b0101101010100101101001010101101001101001100101100110100110010110,
64'b0110100101101001100101101001011000001111111100000000111111110000,
64'b0101101001011010010110100101101001010101010101011010101010101010,
64'b0000000000000000000000000000000011110000000011110000111111110000,
64'b0000000000000000000000000000000010010110100101101001011010010110,
64'b0101010110101010010101011010101000001111111100000000111111110000,
64'b0011110000111100001111000011110011000011110000110011110000111100,
64'b0011001111001100001100111100110000001111111100000000111111110000,
64'b1100001111000011001111000011110011111111111111110000000000000000,
64'b0110100110010110011010011001011011001100001100110011001111001100,
64'b0011001100110011110011001100110000111100110000111100001100111100,
64'b0011001111001100001100111100110010101010101010101010101010101010,
64'b0011001111001100001100111100110010010110100101101001011010010110,
64'b0110011001100110011001100110011000111100110000111100001100111100,
64'b1010101001010101010101011010101000000000111111111111111100000000,
64'b1100001100111100110000110011110011001100110011001100110011001100,
64'b0110100101101001100101101001011010101010010101010101010110101010,
64'b1111000000001111000011111111000001101001100101100110100110010110,
64'b0101101001011010010110100101101000000000111111111111111100000000,
64'b0011110011000011110000110011110000001111111100000000111111110000,
64'b1010010101011010101001010101101001010101101010100101010110101010,
64'b1010010101011010101001010101101000000000111111111111111100000000,
64'b1001011001101001011010011001011000111100001111000011110000111100,
64'b1111000011110000111100001111000000111100110000111100001100111100,
64'b1010010110100101010110100101101001100110100110011001100101100110,
64'b0000111100001111111100001111000010101010101010101010101010101010,
64'b0011110000111100001111000011110011110000111100001111000011110000,
64'b0011001100110011110011001100110010010110100101101001011010010110,
64'b0101101010100101101001010101101000000000000000000000000000000000,
64'b1100001100111100110000110011110001011010010110100101101001011010,
64'b1010101001010101010101011010101001100110011001100110011001100110,
64'b1001100101100110100110010110011010010110100101101001011010010110,
64'b1111000000001111000011111111000010011001011001101001100101100110,
64'b1001100101100110100110010110011010011001011001101001100101100110,
64'b0110011001100110011001100110011011111111000000001111111100000000,
64'b1010010101011010101001010101101000111100110000111100001100111100,
64'b0011001111001100001100111100110010010110011010010110100110010110,
64'b0011001100110011110011001100110001101001100101100110100110010110,
64'b0011110000111100001111000011110000001111111100000000111111110000,
64'b1010010110100101010110100101101011111111111111110000000000000000,
64'b0011001100110011110011001100110000000000111111111111111100000000,
64'b0011110011000011110000110011110001011010010110100101101001011010,
64'b0011001111001100001100111100110001011010101001011010010101011010,
64'b1100001100111100110000110011110011001100001100110011001111001100,
64'b0000000000000000000000000000000010101010010101010101010110101010,
64'b0011001111001100001100111100110011110000111100001111000011110000,
64'b1100001100111100110000110011110001101001100101100110100110010110,
64'b1001011001101001011010011001011011111111111111110000000000000000,
64'b0101010110101010010101011010101011110000000011110000111111110000,
64'b0110100101101001100101101001011010010110011010010110100110010110,
64'b1111000000001111000011111111000010010110011010010110100110010110,
64'b1100110011001100110011001100110000000000111111111111111100000000,
64'b0011001100110011110011001100110000000000000000000000000000000000,
64'b1001100110011001011001100110011001010101010101011010101010101010,
64'b0000000011111111111111110000000010011001011001101001100101100110,
64'b1100110011001100110011001100110011001100001100110011001111001100,
64'b0000000000000000000000000000000010100101101001010101101001011010,
64'b0110100101101001100101101001011010011001100110010110011001100110,
64'b0011110000111100001111000011110001010101101010100101010110101010,
64'b0101101001011010010110100101101011000011001111001100001100111100,
64'b0011110011000011110000110011110000000000000000000000000000000000,
64'b1001100110011001011001100110011010101010010101010101010110101010,
64'b1100001100111100110000110011110010010110011010010110100110010110,
64'b1010101001010101010101011010101010010110011010010110100110010110,
64'b0101101001011010010110100101101001010101010101011010101010101010,
64'b1111000011110000111100001111000010101010101010101010101010101010,
64'b1001011010010110100101101001011011001100110011001100110011001100,
64'b0101010101010101101010101010101001101001011010011001011010010110,
64'b0101101001011010010110100101101000001111000011111111000011110000,
64'b0000000000000000000000000000000010011001011001101001100101100110,
64'b1100001100111100110000110011110010010110100101101001011010010110,
64'b1010010101011010101001010101101010011001100110010110011001100110,
64'b0011001111001100001100111100110000001111111100000000111111110000,
64'b1111000011110000111100001111000010101010010101010101010110101010,
64'b0000111100001111111100001111000010101010101010101010101010101010,
64'b0011110011000011110000110011110011110000000011110000111111110000,
64'b0011001111001100001100111100110010010110100101101001011010010110,
64'b1111000011110000111100001111000000001111111100000000111111110000,
64'b1111111111111111000000000000000001100110100110011001100101100110,
64'b0000000011111111111111110000000000110011001100111100110011001100,
64'b1001011010010110100101101001011010011001011001101001100101100110,
64'b1111000000001111000011111111000000111100110000111100001100111100,
64'b1111000000001111000011111111000010011001011001101001100101100110,
64'b1001100101100110100110010110011010101010010101010101010110101010,
64'b1111111100000000111111110000000000001111000011111111000011110000,
64'b1010010101011010101001010101101000000000000000000000000000000000,
64'b0101010101010101101010101010101010011001100110010110011001100110,
64'b0110011010011001100110010110011001100110011001100110011001100110,
64'b0011110011000011110000110011110000000000111111111111111100000000,
64'b1010010101011010101001010101101001101001100101100110100110010110,
64'b1001011010010110100101101001011000000000111111111111111100000000,
64'b0000000011111111111111110000000011000011110000110011110000111100,
64'b1001011010010110100101101001011001011010010110100101101001011010,
64'b0011001111001100001100111100110001101001011010011001011010010110,
64'b0110100110010110011010011001011011110000000011110000111111110000,
64'b0101101001011010010110100101101001101001011010011001011010010110,
64'b0000000000000000000000000000000000110011001100111100110011001100,
64'b1100110011001100110011001100110001010101101010100101010110101010,
64'b0110011001100110011001100110011010101010101010101010101010101010,
64'b1100110000110011001100111100110010010110100101101001011010010110,
64'b1111000011110000111100001111000010010110100101101001011010010110,
64'b0011110011000011110000110011110011111111111111110000000000000000,
64'b0110011001100110011001100110011010010110011010010110100110010110,
64'b1010101010101010101010101010101011111111111111110000000000000000,
64'b1111111100000000111111110000000010100101010110101010010101011010,
64'b1010101001010101010101011010101010011001011001101001100101100110,
64'b0101010101010101101010101010101011000011001111001100001100111100,
64'b0101010110101010010101011010101010101010010101010101010110101010,
64'b1100001111000011001111000011110001101001100101100110100110010110,
64'b0110100101101001100101101001011001011010010110100101101001011010,
64'b1100001111000011001111000011110010011001100110010110011001100110,
64'b0110100110010110011010011001011011001100110011001100110011001100,
64'b0000111100001111111100001111000001101001100101100110100110010110,
64'b0101010110101010010101011010101011000011001111001100001100111100,
64'b1111000000001111000011111111000000000000000000000000000000000000,
64'b1001011010010110100101101001011010010110011010010110100110010110,
64'b1100110011001100110011001100110010101010101010101010101010101010,
64'b1111111111111111000000000000000001100110100110011001100101100110,
64'b0011001100110011110011001100110011000011110000110011110000111100,
64'b0110011001100110011001100110011011110000000011110000111111110000,
64'b1001100110011001011001100110011000110011001100111100110011001100,
64'b0000111111110000000011111111000010010110011010010110100110010110,
64'b0110100110010110011010011001011000110011110011000011001111001100,
64'b1010010101011010101001010101101000111100001111000011110000111100,
64'b0110100110010110011010011001011001011010010110100101101001011010,
64'b1111111100000000111111110000000000111100110000111100001100111100,
64'b1001100110011001011001100110011011110000000011110000111111110000,
64'b0000000011111111111111110000000000000000000000000000000000000000,
64'b0110100110010110011010011001011000111100110000111100001100111100,
64'b1111000011110000111100001111000001100110011001100110011001100110,
64'b0000000000000000000000000000000011000011110000110011110000111100,
64'b0101101001011010010110100101101010100101010110101010010101011010,
64'b1001011010010110100101101001011010101010010101010101010110101010,
64'b0011110000111100001111000011110001011010010110100101101001011010,
64'b1010101001010101010101011010101010010110011010010110100110010110,
64'b0011110011000011110000110011110010100101101001010101101001011010,
64'b1100110000110011001100111100110000001111111100000000111111110000,
64'b1100001100111100110000110011110000110011110011000011001111001100,
64'b0101010101010101101010101010101011110000000011110000111111110000,
64'b0011110000111100001111000011110010101010010101010101010110101010,
64'b0101010101010101101010101010101010101010101010101010101010101010,
64'b1001011001101001011010011001011011110000000011110000111111110000,
64'b1111111100000000111111110000000010010110100101101001011010010110,
64'b0000000000000000000000000000000000001111111100000000111111110000,
64'b0011001111001100001100111100110001100110100110011001100101100110,
64'b1100001100111100110000110011110000110011001100111100110011001100,
64'b0000111111110000000011111111000010011001011001101001100101100110,
64'b0011001100110011110011001100110000111100110000111100001100111100,
64'b0101101010100101101001010101101010011001011001101001100101100110,
64'b1010010110100101010110100101101010101010010101010101010110101010,
64'b1010010101011010101001010101101011110000111100001111000011110000,
64'b1100110011001100110011001100110010100101010110101010010101011010,
64'b1100110000110011001100111100110011000011110000110011110000111100,
64'b1111000000001111000011111111000001011010101001011010010101011010,
64'b0000111100001111111100001111000011000011001111001100001100111100,
64'b0110100101101001100101101001011011111111111111110000000000000000,
64'b1100110000110011001100111100110010010110011010010110100110010110,
64'b0000111100001111111100001111000000111100110000111100001100111100,
64'b0011110011000011110000110011110011000011001111001100001100111100,
64'b1111000000001111000011111111000001101001011010011001011010010110,
64'b1010010110100101010110100101101011000011110000110011110000111100,
64'b0000111100001111111100001111000001101001011010011001011010010110,
64'b0000000011111111111111110000000010010110100101101001011010010110,
64'b1100110011001100110011001100110010010110100101101001011010010110,
64'b1001011010010110100101101001011011001100001100110011001111001100,
64'b1100001100111100110000110011110000001111111100000000111111110000,
64'b0101101001011010010110100101101001100110100110011001100101100110,
64'b0101101010100101101001010101101001011010101001011010010101011010,
64'b0000000011111111111111110000000000000000000000000000000000000000,
64'b0110100110010110011010011001011010010110011010010110100110010110,
64'b0101101010100101101001010101101001011010101001011010010101011010,
64'b0110011001100110011001100110011001011010101001011010010101011010,
64'b0101101001011010010110100101101011000011001111001100001100111100,
64'b0011110011000011110000110011110010100101010110101010010101011010,
64'b0101101010100101101001010101101001101001100101100110100110010110,
64'b0101010110101010010101011010101001101001100101100110100110010110,
64'b1001011010010110100101101001011011000011001111001100001100111100,
64'b1010010101011010101001010101101000001111000011111111000011110000,
64'b0011110000111100001111000011110010101010010101010101010110101010,
64'b1100001111000011001111000011110011000011110000110011110000111100,
64'b1100001100111100110000110011110001100110100110011001100101100110,
64'b0011110000111100001111000011110010101010101010101010101010101010,
64'b0101101001011010010110100101101000111100110000111100001100111100,
64'b1100001100111100110000110011110001100110100110011001100101100110,
64'b1010101001010101010101011010101001100110100110011001100101100110,
64'b1100001111000011001111000011110001011010101001011010010101011010,
64'b0101010110101010010101011010101011001100001100110011001111001100,
64'b0110100110010110011010011001011000111100110000111100001100111100,
64'b1001100101100110100110010110011000111100110000111100001100111100,
64'b0000111111110000000011111111000000001111111100000000111111110000,
64'b0110011010011001100110010110011001010101101010100101010110101010,
64'b0000111111110000000011111111000010011001100110010110011001100110,
64'b0000111111110000000011111111000010100101010110101010010101011010,
64'b0101101010100101101001010101101001101001011010011001011010010110,
64'b0000111111110000000011111111000001100110011001100110011001100110,
64'b0011001111001100001100111100110011110000000011110000111111110000,
64'b1111000000001111000011111111000001101001011010011001011010010110,
64'b0011001100110011110011001100110001101001011010011001011010010110,
64'b1010010101011010101001010101101001100110100110011001100101100110,
64'b1001100110011001011001100110011010100101101001010101101001011010,
64'b0011110011000011110000110011110001011010101001011010010101011010,
64'b1100001111000011001111000011110001011010101001011010010101011010,
64'b1111111100000000111111110000000001010101101010100101010110101010,
64'b1010010110100101010110100101101000110011001100111100110011001100,
64'b0110011001100110011001100110011000111100001111000011110000111100,
64'b1111000011110000111100001111000001100110100110011001100101100110,
64'b1100001100111100110000110011110011000011001111001100001100111100,
64'b1100001100111100110000110011110010010110100101101001011010010110,
64'b1100001100111100110000110011110000000000111111111111111100000000,
64'b0000111111110000000011111111000001101001100101100110100110010110,
64'b0110011010011001100110010110011001101001100101100110100110010110,
64'b1001011010010110100101101001011001101001011010011001011010010110,
64'b1001100110011001011001100110011010011001011001101001100101100110,
64'b0101010110101010010101011010101001100110100110011001100101100110,
64'b1010010110100101010110100101101001100110100110011001100101100110,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b0101010110101010010101011010101001011010010110100101101001011010,
64'b0101101010100101101001010101101010100101010110101010010101011010,
64'b0000111100001111111100001111000011000011110000110011110000111100,
64'b1111111100000000111111110000000001011010101001011010010101011010,
64'b1001100101100110100110010110011011000011001111001100001100111100,
64'b0011110000111100001111000011110011111111111111110000000000000000,
64'b0000111111110000000011111111000010010110011010010110100110010110,
64'b1111111100000000111111110000000000111100110000111100001100111100,
64'b1001100110011001011001100110011011000011001111001100001100111100,
64'b1001100110011001011001100110011001101001011010011001011010010110,
64'b1001011010010110100101101001011011000011110000110011110000111100,
64'b0011001100110011110011001100110001101001011010011001011010010110,
64'b0101101001011010010110100101101010010110100101101001011010010110,
64'b1001100110011001011001100110011001010101101010100101010110101010,
64'b1100110000110011001100111100110000000000000000000000000000000000,
64'b0101010110101010010101011010101011111111111111110000000000000000,
64'b0101010101010101101010101010101001101001100101100110100110010110,
64'b1100001111000011001111000011110000110011110011000011001111001100,
64'b0000111111110000000011111111000011001100001100110011001111001100,
64'b0000000011111111111111110000000010011001011001101001100101100110,
64'b1111111111111111000000000000000001100110011001100110011001100110,
64'b0011110000111100001111000011110010101010101010101010101010101010,
64'b1001011010010110100101101001011001100110100110011001100101100110,
64'b0110100110010110011010011001011010101010010101010101010110101010,
64'b1111000011110000111100001111000001101001011010011001011010010110,
64'b1001100101100110100110010110011010100101010110101010010101011010,
64'b0101101001011010010110100101101001010101010101011010101010101010,
64'b0110100110010110011010011001011011001100001100110011001111001100,
64'b0110100110010110011010011001011011110000000011110000111111110000,
64'b1100001111000011001111000011110010011001011001101001100101100110,
64'b1100110000110011001100111100110001100110011001100110011001100110,
64'b0110011001100110011001100110011011000011001111001100001100111100,
64'b1111000011110000111100001111000001100110011001100110011001100110,
64'b1001011001101001011010011001011000000000111111111111111100000000,
64'b0101010101010101101010101010101000111100110000111100001100111100,
64'b0110011010011001100110010110011001100110011001100110011001100110,
64'b0011001111001100001100111100110010010110100101101001011010010110,
64'b1111111111111111000000000000000001101001011010011001011010010110,
64'b1111000011110000111100001111000001010101101010100101010110101010,
64'b0101010110101010010101011010101001100110011001100110011001100110,
64'b1111000011110000111100001111000010100101101001010101101001011010,
64'b1100110011001100110011001100110010101010010101010101010110101010,
64'b0000000011111111111111110000000001101001011010011001011010010110,
64'b1100110011001100110011001100110000111100001111000011110000111100,
64'b0101101010100101101001010101101011110000000011110000111111110000,
64'b1111000000001111000011111111000000111100001111000011110000111100,
64'b0000000000000000000000000000000011111111111111110000000000000000,
64'b1001011001101001011010011001011001011010101001011010010101011010,
64'b1100110011001100110011001100110010010110100101101001011010010110,
64'b1010101010101010101010101010101011000011001111001100001100111100,
64'b0000000011111111111111110000000011000011001111001100001100111100,
64'b1001100101100110100110010110011001100110011001100110011001100110,
64'b0011001100110011110011001100110010010110100101101001011010010110,
64'b1111111100000000111111110000000000110011110011000011001111001100,
64'b1111000011110000111100001111000010011001100110010110011001100110,
64'b1111111111111111000000000000000001101001100101100110100110010110,
64'b0101101001011010010110100101101010100101010110101010010101011010,
64'b1100110000110011001100111100110000000000111111111111111100000000,
64'b1010101001010101010101011010101010100101010110101010010101011010,
64'b1010101010101010101010101010101000000000000000000000000000000000,
64'b0011110011000011110000110011110001100110100110011001100101100110,
64'b0101101001011010010110100101101001101001100101100110100110010110,
64'b1100110011001100110011001100110011110000000011110000111111110000,
64'b1111111111111111000000000000000011110000000011110000111111110000,
64'b1001011010010110100101101001011000111100001111000011110000111100,
64'b1001011010010110100101101001011010100101010110101010010101011010,
64'b1001100101100110100110010110011011000011001111001100001100111100,
64'b0000111100001111111100001111000011001100001100110011001111001100,
64'b0000111100001111111100001111000010011001011001101001100101100110,
64'b1111000000001111000011111111000010100101010110101010010101011010,
64'b1100001100111100110000110011110000110011110011000011001111001100,
64'b1001011010010110100101101001011001101001100101100110100110010110,
64'b0101101010100101101001010101101000111100110000111100001100111100,
64'b0000000000000000000000000000000000110011110011000011001111001100,
64'b0011110011000011110000110011110000110011110011000011001111001100,
64'b1111111111111111000000000000000000001111111100000000111111110000,
64'b0000000011111111111111110000000010101010101010101010101010101010,
64'b1010010101011010101001010101101001101001100101100110100110010110,
64'b1010010101011010101001010101101011001100001100110011001111001100,
64'b0000111111110000000011111111000011110000000011110000111111110000,
64'b0000111100001111111100001111000000001111000011111111000011110000,
64'b0101101010100101101001010101101001101001011010011001011010010110,
64'b1100001100111100110000110011110011001100001100110011001111001100,
64'b1001011010010110100101101001011000001111000011111111000011110000,
64'b1100110000110011001100111100110000111100110000111100001100111100,
64'b1111000011110000111100001111000011110000000011110000111111110000,
64'b0101101010100101101001010101101010100101101001010101101001011010,
64'b0101010110101010010101011010101000001111000011111111000011110000,
64'b1010010110100101010110100101101000000000111111111111111100000000,
64'b0101010110101010010101011010101011001100110011001100110011001100,
64'b0101010110101010010101011010101011000011001111001100001100111100,
64'b0000000011111111111111110000000000001111000011111111000011110000,
64'b1100110011001100110011001100110010101010010101010101010110101010,
64'b0000111100001111111100001111000001010101101010100101010110101010,
64'b0110100110010110011010011001011001101001100101100110100110010110,
64'b0011001111001100001100111100110010100101101001010101101001011010,
64'b0000111100001111111100001111000001010101101010100101010110101010,
64'b0000000000000000000000000000000001011010101001011010010101011010,
64'b0110100101101001100101101001011010101010010101010101010110101010,
64'b0011110000111100001111000011110010011001011001101001100101100110,
64'b0011110000111100001111000011110001010101101010100101010110101010,
64'b0011110011000011110000110011110001010101010101011010101010101010,
64'b1001100101100110100110010110011001011010010110100101101001011010,
64'b0000000000000000000000000000000000001111111100000000111111110000,
64'b0101010101010101101010101010101011111111000000001111111100000000,
64'b0101101001011010010110100101101010011001100110010110011001100110,
64'b1111111100000000111111110000000010011001100110010110011001100110,
64'b1001011001101001011010011001011000111100110000111100001100111100,
64'b0000111100001111111100001111000000110011110011000011001111001100,
64'b1111111100000000111111110000000010011001100110010110011001100110,
64'b1010101010101010101010101010101011001100001100110011001111001100,
64'b1100001100111100110000110011110010011001100110010110011001100110,
64'b1010010101011010101001010101101001101001011010011001011010010110,
64'b0000111111110000000011111111000000110011001100111100110011001100,
64'b1111000000001111000011111111000011001100110011001100110011001100,
64'b0110100101101001100101101001011010011001011001101001100101100110,
64'b0000000000000000000000000000000011111111000000001111111100000000,
64'b0110011001100110011001100110011011111111111111110000000000000000,
64'b1001100101100110100110010110011000111100001111000011110000111100,
64'b1111111111111111000000000000000010010110100101101001011010010110,
64'b0011110011000011110000110011110001011010101001011010010101011010,
64'b0101010110101010010101011010101010100101101001010101101001011010,
64'b0101010101010101101010101010101000111100001111000011110000111100,
64'b1100110011001100110011001100110010100101101001010101101001011010,
64'b1111000000001111000011111111000010010110100101101001011010010110,
64'b1100110000110011001100111100110001101001100101100110100110010110,
64'b0000000011111111111111110000000001011010010110100101101001011010,
64'b0000000011111111111111110000000001011010010110100101101001011010,
64'b0110100110010110011010011001011011000011110000110011110000111100,
64'b1010101010101010101010101010101000000000000000000000000000000000,
64'b1001011010010110100101101001011010101010101010101010101010101010,
64'b1100001111000011001111000011110010100101010110101010010101011010,
64'b0000000000000000000000000000000011000011001111001100001100111100,
64'b0101101010100101101001010101101011001100001100110011001111001100,
64'b1001100110011001011001100110011010011001011001101001100101100110,
64'b1100110011001100110011001100110010100101010110101010010101011010,
64'b0101101001011010010110100101101000110011110011000011001111001100,
64'b0000000011111111111111110000000001101001100101100110100110010110,
64'b1010010110100101010110100101101000111100110000111100001100111100,
64'b0101010101010101101010101010101000110011110011000011001111001100,
64'b0101010101010101101010101010101000110011110011000011001111001100,
64'b1001011001101001011010011001011000001111111100000000111111110000,
64'b1100110011001100110011001100110010101010101010101010101010101010,
64'b1111000000001111000011111111000000001111111100000000111111110000,
64'b1010101010101010101010101010101011000011001111001100001100111100,
64'b0101101010100101101001010101101011001100001100110011001111001100,
64'b1001100110011001011001100110011000001111111100000000111111110000,
64'b0000000011111111111111110000000000000000111111111111111100000000,
64'b1001011001101001011010011001011011000011110000110011110000111100,
64'b1100110011001100110011001100110010101010101010101010101010101010,
64'b0101101001011010010110100101101000111100110000111100001100111100,
64'b0000111100001111111100001111000010101010101010101010101010101010,
64'b0000111111110000000011111111000001010101010101011010101010101010,
64'b0110011010011001100110010110011011001100110011001100110011001100,
64'b0110100110010110011010011001011001101001100101100110100110010110,
64'b1001100101100110100110010110011010010110100101101001011010010110,
64'b1111000011110000111100001111000000000000111111111111111100000000,
64'b1100110011001100110011001100110011110000000011110000111111110000,
64'b1001011010010110100101101001011000001111000011111111000011110000,
64'b0000111100001111111100001111000010101010010101010101010110101010,
64'b0101010110101010010101011010101011111111111111110000000000000000,
64'b0000000000000000000000000000000010100101010110101010010101011010,
64'b1001011010010110100101101001011001100110011001100110011001100110,
64'b0110100110010110011010011001011011110000000011110000111111110000,
64'b1111000000001111000011111111000001100110011001100110011001100110,
64'b1010010110100101010110100101101011001100110011001100110011001100,
64'b1010010101011010101001010101101001011010010110100101101001011010,
64'b1111111111111111000000000000000000111100110000111100001100111100,
64'b1010010101011010101001010101101011000011001111001100001100111100,
64'b0000111100001111111100001111000001010101010101011010101010101010,
64'b0101101001011010010110100101101010101010010101010101010110101010,
64'b1001100110011001011001100110011001010101101010100101010110101010,
64'b0110011010011001100110010110011010011001100110010110011001100110,
64'b1001100101100110100110010110011010101010101010101010101010101010,
64'b1001011001101001011010011001011001100110100110011001100101100110,
64'b0000111111110000000011111111000000111100001111000011110000111100,
64'b0110011010011001100110010110011000000000111111111111111100000000,
64'b0000111111110000000011111111000010010110100101101001011010010110,
64'b1001011010010110100101101001011011110000111100001111000011110000,
64'b0000000000000000000000000000000000110011110011000011001111001100,
64'b0110100110010110011010011001011011110000000011110000111111110000,
64'b0000000000000000000000000000000010100101010110101010010101011010,
64'b0101010110101010010101011010101001100110011001100110011001100110,
64'b1001100101100110100110010110011010011001100110010110011001100110,
64'b0011110000111100001111000011110010011001100110010110011001100110,
64'b0110100101101001100101101001011000111100001111000011110000111100,
64'b0110100101101001100101101001011001100110011001100110011001100110,
64'b0011110011000011110000110011110011000011110000110011110000111100,
64'b1010101001010101010101011010101010100101010110101010010101011010,
64'b1100001111000011001111000011110011111111111111110000000000000000,
64'b1010101001010101010101011010101001101001100101100110100110010110,
64'b1100001100111100110000110011110011111111000000001111111100000000,
64'b0000000000000000000000000000000000001111000011111111000011110000,
64'b0011110011000011110000110011110000000000111111111111111100000000,
64'b0000000000000000000000000000000010011001011001101001100101100110,
64'b0110100110010110011010011001011010010110100101101001011010010110,
64'b0110100101101001100101101001011000111100001111000011110000111100,
64'b0101010101010101101010101010101010010110100101101001011010010110,
64'b0101101010100101101001010101101010100101010110101010010101011010,
64'b0110100101101001100101101001011000111100001111000011110000111100,
64'b1100110011001100110011001100110000001111111100000000111111110000,
64'b0101010101010101101010101010101001100110100110011001100101100110,
64'b1111111100000000111111110000000000000000000000000000000000000000,
64'b1001011010010110100101101001011010010110011010010110100110010110,
64'b0101010101010101101010101010101011111111111111110000000000000000,
64'b0110011010011001100110010110011011111111000000001111111100000000,
64'b1001100110011001011001100110011001010101010101011010101010101010,
64'b0011001111001100001100111100110010010110100101101001011010010110,
64'b1100110011001100110011001100110011000011001111001100001100111100,
64'b0110100110010110011010011001011000001111111100000000111111110000,
64'b0011110011000011110000110011110011000011001111001100001100111100,
64'b1111111100000000111111110000000011001100001100110011001111001100,
64'b0110100101101001100101101001011000001111111100000000111111110000,
64'b1100110000110011001100111100110000000000111111111111111100000000,
64'b0000000000000000000000000000000011000011110000110011110000111100,
64'b0000111100001111111100001111000010101010101010101010101010101010,
64'b1100110000110011001100111100110000111100110000111100001100111100,
64'b1100001100111100110000110011110010101010101010101010101010101010,
64'b0000111111110000000011111111000001010101010101011010101010101010,
64'b1111111100000000111111110000000011001100110011001100110011001100,
64'b1100001100111100110000110011110001101001100101100110100110010110,
64'b1111000011110000111100001111000000000000000000000000000000000000,
64'b0011110011000011110000110011110010101010010101010101010110101010,
64'b1111000000001111000011111111000010101010101010101010101010101010,
64'b0101010101010101101010101010101010010110100101101001011010010110,
64'b1100001100111100110000110011110010101010101010101010101010101010,
64'b1010010110100101010110100101101001101001100101100110100110010110,
64'b1010101010101010101010101010101001101001100101100110100110010110,
64'b1111111100000000111111110000000000111100001111000011110000111100,
64'b1010010110100101010110100101101011111111000000001111111100000000,
64'b0101101010100101101001010101101001101001100101100110100110010110,
64'b0000000011111111111111110000000010101010010101010101010110101010,
64'b1111111111111111000000000000000000110011110011000011001111001100,
64'b0000111111110000000011111111000001011010010110100101101001011010,
64'b1010010110100101010110100101101001011010101001011010010101011010,
64'b0101101010100101101001010101101010011001100110010110011001100110,
64'b1111000011110000111100001111000000111100110000111100001100111100,
64'b1111111111111111000000000000000001011010101001011010010101011010,
64'b0101101001011010010110100101101011001100001100110011001111001100,
64'b1010010110100101010110100101101010101010101010101010101010101010,
64'b1010101010101010101010101010101011110000000011110000111111110000,
64'b1010010110100101010110100101101001010101101010100101010110101010,
64'b0011110011000011110000110011110011110000111100001111000011110000,
64'b0110100101101001100101101001011000110011001100111100110011001100,
64'b0011001111001100001100111100110001010101101010100101010110101010,
64'b1100001100111100110000110011110011001100001100110011001111001100,
64'b1100110011001100110011001100110010101010101010101010101010101010,
64'b1100001111000011001111000011110001100110100110011001100101100110,
64'b1100110000110011001100111100110010010110100101101001011010010110,
64'b0000111100001111111100001111000001011010101001011010010101011010,
64'b1001100110011001011001100110011001100110100110011001100101100110,
64'b1001100110011001011001100110011010100101101001010101101001011010,
64'b1010010110100101010110100101101001100110011001100110011001100110,
64'b1010101010101010101010101010101000000000111111111111111100000000,
64'b0110100110010110011010011001011010011001100110010110011001100110,
64'b0101010110101010010101011010101011111111000000001111111100000000,
64'b0110011001100110011001100110011011110000111100001111000011110000,
64'b1100001100111100110000110011110010011001100110010110011001100110,
64'b1001100110011001011001100110011000001111000011111111000011110000,
64'b0110100110010110011010011001011001100110011001100110011001100110,
64'b1010010101011010101001010101101011000011110000110011110000111100,
64'b1010010110100101010110100101101001101001100101100110100110010110,
64'b0101010110101010010101011010101011001100001100110011001111001100,
64'b1001011010010110100101101001011001101001011010011001011010010110,
64'b1001011010010110100101101001011010011001011001101001100101100110,
64'b1001100101100110100110010110011010010110100101101001011010010110,
64'b0110011001100110011001100110011011111111111111110000000000000000,
64'b0011110011000011110000110011110010010110100101101001011010010110,
64'b0011001100110011110011001100110001010101010101011010101010101010,
64'b0011110000111100001111000011110011111111000000001111111100000000,
64'b1111000000001111000011111111000000111100001111000011110000111100,
64'b0011110000111100001111000011110001010101101010100101010110101010,
64'b0110100110010110011010011001011010010110100101101001011010010110,
64'b0011110000111100001111000011110011111111111111110000000000000000,
64'b1001100101100110100110010110011000111100110000111100001100111100,
64'b1100001100111100110000110011110001010101101010100101010110101010,
64'b0101101010100101101001010101101011110000000011110000111111110000,
64'b1100001111000011001111000011110001101001100101100110100110010110,
64'b0101010110101010010101011010101001010101010101011010101010101010,
64'b1111000011110000111100001111000011001100110011001100110011001100,
64'b1010101001010101010101011010101000110011110011000011001111001100,
64'b0101010101010101101010101010101011000011110000110011110000111100,
64'b1010101010101010101010101010101001011010101001011010010101011010,
64'b0110011001100110011001100110011001101001011010011001011010010110,
64'b1100110011001100110011001100110001011010101001011010010101011010,
64'b0101101001011010010110100101101001011010010110100101101001011010,
64'b0101010101010101101010101010101010101010101010101010101010101010,
64'b0110100101101001100101101001011001011010101001011010010101011010,
64'b1010101010101010101010101010101010011001100110010110011001100110,
64'b0101010110101010010101011010101000000000111111111111111100000000,
64'b1010010110100101010110100101101010010110011010010110100110010110,
64'b0000111111110000000011111111000011001100110011001100110011001100,
64'b0011001111001100001100111100110001011010010110100101101001011010,
64'b0110100101101001100101101001011000001111000011111111000011110000,
64'b0110100101101001100101101001011000001111111100000000111111110000,
64'b0110100110010110011010011001011001100110100110011001100101100110,
64'b0101101010100101101001010101101001101001100101100110100110010110,
64'b1001100101100110100110010110011001100110100110011001100101100110,
64'b1010101010101010101010101010101010011001011001101001100101100110,
64'b1001011001101001011010011001011001100110011001100110011001100110,
64'b1100001100111100110000110011110011001100001100110011001111001100,
64'b0011110011000011110000110011110010010110100101101001011010010110,
64'b1010101010101010101010101010101001010101010101011010101010101010,
64'b0011001100110011110011001100110010010110011010010110100110010110,
64'b0011110000111100001111000011110001011010010110100101101001011010,
64'b1100001111000011001111000011110000110011110011000011001111001100,
64'b1001100101100110100110010110011011111111000000001111111100000000,
64'b0110011010011001100110010110011010101010010101010101010110101010,
64'b1001100110011001011001100110011011000011110000110011110000111100,
64'b1010101010101010101010101010101010010110011010010110100110010110,
64'b0000000011111111111111110000000011000011110000110011110000111100,
64'b0101010110101010010101011010101010010110100101101001011010010110,
64'b0011110011000011110000110011110010010110100101101001011010010110,
64'b0101101010100101101001010101101000001111000011111111000011110000,
64'b1111000000001111000011111111000001101001100101100110100110010110,
64'b0110011001100110011001100110011011001100110011001100110011001100,
64'b1111000011110000111100001111000010010110011010010110100110010110,
64'b1010010101011010101001010101101010011001011001101001100101100110,
64'b0000111111110000000011111111000000001111000011111111000011110000,
64'b0110100101101001100101101001011011111111111111110000000000000000,
64'b1100001111000011001111000011110000110011001100111100110011001100,
64'b1001011010010110100101101001011010100101010110101010010101011010,
64'b0110011001100110011001100110011010010110011010010110100110010110,
64'b1111111111111111000000000000000010100101010110101010010101011010,
64'b0110011001100110011001100110011001101001100101100110100110010110,
64'b1111000000001111000011111111000001101001100101100110100110010110,
64'b0110011010011001100110010110011011111111000000001111111100000000,
64'b1010101001010101010101011010101010010110011010010110100110010110,
64'b1001011010010110100101101001011011110000111100001111000011110000,
64'b1111111100000000111111110000000000111100110000111100001100111100,
64'b1100110000110011001100111100110001101001011010011001011010010110,
64'b0000000011111111111111110000000011111111000000001111111100000000,
64'b1100001100111100110000110011110010101010101010101010101010101010,
64'b1010010101011010101001010101101001011010010110100101101001011010,
64'b0110100110010110011010011001011001100110100110011001100101100110,
64'b0011110000111100001111000011110000111100110000111100001100111100,
64'b0000000000000000000000000000000001100110100110011001100101100110,
64'b1001011010010110100101101001011011000011001111001100001100111100,
64'b0000000011111111111111110000000000111100110000111100001100111100,
64'b0110100101101001100101101001011011111111111111110000000000000000,
64'b1001100110011001011001100110011000111100110000111100001100111100,
64'b0110100110010110011010011001011001010101101010100101010110101010,
64'b1111111111111111000000000000000011110000000011110000111111110000,
64'b0000111100001111111100001111000001101001100101100110100110010110,
64'b0101010101010101101010101010101001010101010101011010101010101010,
64'b0101101010100101101001010101101011001100110011001100110011001100,
64'b1100110000110011001100111100110000110011110011000011001111001100,
64'b0011110011000011110000110011110011000011110000110011110000111100,
64'b0000111111110000000011111111000001011010101001011010010101011010,
64'b0000000000000000000000000000000001101001011010011001011010010110,
64'b1100001100111100110000110011110010100101010110101010010101011010,
64'b0110100101101001100101101001011011000011001111001100001100111100,
64'b0011110011000011110000110011110000110011001100111100110011001100,
64'b1111000000001111000011111111000010010110011010010110100110010110,
64'b0000111100001111111100001111000001100110011001100110011001100110,
64'b1001011001101001011010011001011001101001011010011001011010010110,
64'b1100001100111100110000110011110001101001011010011001011010010110,
64'b0011001111001100001100111100110000000000000000000000000000000000,
64'b1001100110011001011001100110011001011010010110100101101001011010,
64'b1100001111000011001111000011110000001111111100000000111111110000,
64'b1100001111000011001111000011110001100110100110011001100101100110,
64'b1100110000110011001100111100110010010110011010010110100110010110,
64'b1111111111111111000000000000000010011001011001101001100101100110,
64'b0000000000000000000000000000000010100101010110101010010101011010,
64'b0000000011111111111111110000000011110000000011110000111111110000,
64'b0110011001100110011001100110011011110000111100001111000011110000,
64'b0101101001011010010110100101101010010110011010010110100110010110,
64'b0101101010100101101001010101101010010110100101101001011010010110,
64'b0000000000000000000000000000000011000011001111001100001100111100,
64'b1001100110011001011001100110011001101001100101100110100110010110,
64'b0011110011000011110000110011110010101010101010101010101010101010,
64'b1010010110100101010110100101101000110011110011000011001111001100,
64'b0110011010011001100110010110011000000000111111111111111100000000,
64'b0110011010011001100110010110011011000011110000110011110000111100,
64'b0110100110010110011010011001011010010110011010010110100110010110,
64'b0101010101010101101010101010101001101001011010011001011010010110,
64'b1010101010101010101010101010101000110011110011000011001111001100,
64'b0011110000111100001111000011110010101010010101010101010110101010,
64'b1010101001010101010101011010101001010101101010100101010110101010,
64'b1100001111000011001111000011110000111100110000111100001100111100,
64'b1100001100111100110000110011110001101001100101100110100110010110,
64'b0011110011000011110000110011110011110000000011110000111111110000,
64'b1111111100000000111111110000000000111100110000111100001100111100,
64'b0110100101101001100101101001011011001100110011001100110011001100,
64'b0000000011111111111111110000000000001111000011111111000011110000,
64'b1010101010101010101010101010101011111111111111110000000000000000,
64'b1010101010101010101010101010101010100101010110101010010101011010,
64'b0101101001011010010110100101101010010110011010010110100110010110,
64'b0011001100110011110011001100110001101001100101100110100110010110,
64'b0110011001100110011001100110011001011010010110100101101001011010,
64'b0000111111110000000011111111000010011001100110010110011001100110,
64'b0011001100110011110011001100110010011001100110010110011001100110,
64'b1010010101011010101001010101101011110000000011110000111111110000,
64'b0101101010100101101001010101101010010110011010010110100110010110,
64'b1111000000001111000011111111000000000000111111111111111100000000,
64'b0101010101010101101010101010101001011010101001011010010101011010,
64'b1100001100111100110000110011110001011010010110100101101001011010,
64'b0101010101010101101010101010101011111111000000001111111100000000,
64'b0110011001100110011001100110011010101010101010101010101010101010,
64'b1100110011001100110011001100110001100110100110011001100101100110,
64'b0011001111001100001100111100110000111100110000111100001100111100,
64'b1111000011110000111100001111000010010110011010010110100110010110,
64'b1001011010010110100101101001011000110011110011000011001111001100,
64'b0110100110010110011010011001011010010110100101101001011010010110,
64'b1100110000110011001100111100110010010110100101101001011010010110,
64'b1001011010010110100101101001011010101010010101010101010110101010,
64'b1100001100111100110000110011110010010110011010010110100110010110,
64'b0011110000111100001111000011110001010101010101011010101010101010,
64'b1010010101011010101001010101101001100110100110011001100101100110,
64'b0110100101101001100101101001011010011001011001101001100101100110,
64'b0101010101010101101010101010101011111111111111110000000000000000,
64'b0101010101010101101010101010101011001100110011001100110011001100,
64'b0011001100110011110011001100110011000011110000110011110000111100,
64'b1100001100111100110000110011110001011010101001011010010101011010,
64'b0000000011111111111111110000000010010110011010010110100110010110,
64'b1100001100111100110000110011110001011010010110100101101001011010,
64'b1111111100000000111111110000000011000011001111001100001100111100,
64'b0011001111001100001100111100110011000011001111001100001100111100,
64'b1001100110011001011001100110011000110011001100111100110011001100,
64'b1111111100000000111111110000000010010110011010010110100110010110,
64'b1001100110011001011001100110011001100110011001100110011001100110,
64'b0000111100001111111100001111000001101001011010011001011010010110,
64'b1111000011110000111100001111000001101001011010011001011010010110,
64'b1111111111111111000000000000000000000000000000000000000000000000,
64'b1010010110100101010110100101101001011010010110100101101001011010,
64'b1001100110011001011001100110011000001111111100000000111111110000,
64'b1001011010010110100101101001011001100110100110011001100101100110,
64'b0000000000000000000000000000000010010110011010010110100110010110,
64'b1010010101011010101001010101101010011001011001101001100101100110,
64'b0101010101010101101010101010101000110011110011000011001111001100,
64'b0000111100001111111100001111000011001100110011001100110011001100,
64'b0011110000111100001111000011110000000000111111111111111100000000,
64'b0101010101010101101010101010101010011001011001101001100101100110,
64'b0011110000111100001111000011110000000000111111111111111100000000,
64'b0101010110101010010101011010101000000000000000000000000000000000,
64'b0101010110101010010101011010101001011010010110100101101001011010,
64'b0000000000000000000000000000000000110011001100111100110011001100,
64'b1001100101100110100110010110011011110000000011110000111111110000,
64'b1001011010010110100101101001011011000011001111001100001100111100,
64'b0110100110010110011010011001011000001111111100000000111111110000,
64'b0000000000000000000000000000000001101001100101100110100110010110,
64'b0011001111001100001100111100110010010110100101101001011010010110,
64'b0000111100001111111100001111000001100110011001100110011001100110,
64'b0110100101101001100101101001011011001100001100110011001111001100,
64'b0101010101010101101010101010101000001111111100000000111111110000,
64'b1100001111000011001111000011110001100110011001100110011001100110,
64'b0011001100110011110011001100110001101001100101100110100110010110,
64'b1111000000001111000011111111000001101001100101100110100110010110,
64'b0000000011111111111111110000000000000000000000000000000000000000,
64'b1001100110011001011001100110011001101001011010011001011010010110,
64'b0000000000000000000000000000000001101001100101100110100110010110,
64'b0000000011111111111111110000000010011001011001101001100101100110,
64'b1111000011110000111100001111000011001100110011001100110011001100,
64'b1111111111111111000000000000000011000011001111001100001100111100,
64'b1111000011110000111100001111000011000011001111001100001100111100,
64'b1001011001101001011010011001011000111100001111000011110000111100,
64'b0101010101010101101010101010101000001111000011111111000011110000,
64'b1001011001101001011010011001011010101010010101010101010110101010,
64'b1010101001010101010101011010101000111100001111000011110000111100,
64'b1100110000110011001100111100110000111100110000111100001100111100,
64'b0110100101101001100101101001011000111100110000111100001100111100,
64'b0110011010011001100110010110011000000000000000000000000000000000,
64'b0000111100001111111100001111000011000011001111001100001100111100,
64'b0110100101101001100101101001011010010110011010010110100110010110,
64'b0011110000111100001111000011110011000011110000110011110000111100,
64'b1001100110011001011001100110011011110000111100001111000011110000,
64'b1111111111111111000000000000000011110000000011110000111111110000,
64'b0101010110101010010101011010101000001111111100000000111111110000,
64'b1001011001101001011010011001011000001111111100000000111111110000,
64'b0110011001100110011001100110011011111111000000001111111100000000,
64'b1001011001101001011010011001011010011001100110010110011001100110,
64'b1001100110011001011001100110011010100101010110101010010101011010,
64'b1010010110100101010110100101101011110000000011110000111111110000,
64'b0110100110010110011010011001011001011010101001011010010101011010,
64'b0110100101101001100101101001011010101010101010101010101010101010,
64'b0101010110101010010101011010101011110000000011110000111111110000,
64'b0110100110010110011010011001011000111100110000111100001100111100,
64'b1010010101011010101001010101101010100101010110101010010101011010,
64'b0011110000111100001111000011110001010101101010100101010110101010,
64'b1010101010101010101010101010101000000000111111111111111100000000,
64'b0110011001100110011001100110011001010101101010100101010110101010,
64'b1111111100000000111111110000000001101001100101100110100110010110,
64'b1010101001010101010101011010101011000011001111001100001100111100,
64'b1100110011001100110011001100110011001100001100110011001111001100,
64'b1001100110011001011001100110011001101001100101100110100110010110,
64'b0000111100001111111100001111000010010110100101101001011010010110,
64'b0101010101010101101010101010101010100101101001010101101001011010,
64'b1111000011110000111100001111000001010101101010100101010110101010,
64'b0000000000000000000000000000000010011001011001101001100101100110,
64'b1111111100000000111111110000000010011001011001101001100101100110,
64'b0000111111110000000011111111000010100101010110101010010101011010,
64'b1100001111000011001111000011110011111111000000001111111100000000,
64'b0011001100110011110011001100110000000000000000000000000000000000,
64'b0011110000111100001111000011110001100110011001100110011001100110,
64'b1001011010010110100101101001011000111100110000111100001100111100,
64'b0000111111110000000011111111000011110000000011110000111111110000,
64'b1010101001010101010101011010101000001111000011111111000011110000,
64'b0011001100110011110011001100110010010110011010010110100110010110,
64'b1100001111000011001111000011110011000011001111001100001100111100,
64'b1010010101011010101001010101101000110011110011000011001111001100,
64'b0110011001100110011001100110011010011001100110010110011001100110,
64'b1001100110011001011001100110011011000011110000110011110000111100,
64'b0011110000111100001111000011110011000011110000110011110000111100,
64'b1100001100111100110000110011110011001100001100110011001111001100,
64'b1100001111000011001111000011110011111111111111110000000000000000,
64'b1010010110100101010110100101101000000000000000000000000000000000,
64'b1010010101011010101001010101101000111100001111000011110000111100,
64'b1010101001010101010101011010101001011010101001011010010101011010,
64'b0011110000111100001111000011110010101010010101010101010110101010,
64'b1100001100111100110000110011110001010101101010100101010110101010,
64'b0101010101010101101010101010101010010110011010010110100110010110,
64'b0011001100110011110011001100110001011010101001011010010101011010,
64'b1010010110100101010110100101101000001111000011111111000011110000,
64'b0000111111110000000011111111000000111100001111000011110000111100,
64'b1010010110100101010110100101101010100101010110101010010101011010,
64'b0110011010011001100110010110011010100101010110101010010101011010,
64'b0011001111001100001100111100110010100101101001010101101001011010,
64'b1100001111000011001111000011110010101010101010101010101010101010,
64'b0110011010011001100110010110011010101010101010101010101010101010,
64'b1001100101100110100110010110011000001111111100000000111111110000,
64'b1001100110011001011001100110011011001100001100110011001111001100,
64'b1010010101011010101001010101101010011001100110010110011001100110,
64'b1111000000001111000011111111000010011001100110010110011001100110,
64'b1100110011001100110011001100110000111100110000111100001100111100,
64'b0101101001011010010110100101101001100110100110011001100101100110,
64'b1001100101100110100110010110011001010101101010100101010110101010,
64'b1010101001010101010101011010101010100101010110101010010101011010,
64'b0011001111001100001100111100110011001100001100110011001111001100,
64'b0110100101101001100101101001011011001100001100110011001111001100,
64'b1010010110100101010110100101101000110011110011000011001111001100,
64'b0000111111110000000011111111000001100110011001100110011001100110,
64'b0110100101101001100101101001011011001100110011001100110011001100,
64'b1001011010010110100101101001011011111111000000001111111100000000,
64'b0011110000111100001111000011110010100101101001010101101001011010,
64'b0110011010011001100110010110011010010110100101101001011010010110,
64'b0000000011111111111111110000000010010110100101101001011010010110,
64'b0101101001011010010110100101101001011010101001011010010101011010,
64'b0011001111001100001100111100110001101001011010011001011010010110,
64'b1100001111000011001111000011110010011001100110010110011001100110,
64'b0011001100110011110011001100110011001100001100110011001111001100,
64'b1010010110100101010110100101101000001111000011111111000011110000,
64'b1100001100111100110000110011110010100101101001010101101001011010,
64'b1001100101100110100110010110011010100101101001010101101001011010,
64'b1010101001010101010101011010101000111100001111000011110000111100,
64'b1100001100111100110000110011110011110000111100001111000011110000,
64'b0110100110010110011010011001011000000000000000000000000000000000,
64'b0000111111110000000011111111000010011001011001101001100101100110,
64'b1100001111000011001111000011110001101001100101100110100110010110,
64'b0101010101010101101010101010101011000011001111001100001100111100,
64'b1001100101100110100110010110011011001100001100110011001111001100,
64'b0000111100001111111100001111000001101001100101100110100110010110,
64'b0000111111110000000011111111000010010110100101101001011010010110,
64'b0101101001011010010110100101101010100101101001010101101001011010,
64'b1001100101100110100110010110011001010101101010100101010110101010,
64'b0101101010100101101001010101101010011001011001101001100101100110,
64'b1100001111000011001111000011110010011001011001101001100101100110,
64'b0011001100110011110011001100110010100101010110101010010101011010,
64'b0101101010100101101001010101101011111111000000001111111100000000,
64'b1100001100111100110000110011110000000000000000000000000000000000,
64'b0000111111110000000011111111000001101001011010011001011010010110,
64'b1100001111000011001111000011110011111111111111110000000000000000,
64'b1001100110011001011001100110011000001111111100000000111111110000,
64'b0101101001011010010110100101101001010101101010100101010110101010,
64'b0000000000000000000000000000000001010101010101011010101010101010,
64'b0011110011000011110000110011110010100101010110101010010101011010,
64'b1100001100111100110000110011110010010110011010010110100110010110,
64'b1100001100111100110000110011110000111100001111000011110000111100,
64'b1100001100111100110000110011110011110000111100001111000011110000,
64'b1001100101100110100110010110011010011001011001101001100101100110,
64'b1100110011001100110011001100110000111100001111000011110000111100,
64'b1100110011001100110011001100110000001111111100000000111111110000,
64'b1010101010101010101010101010101011001100110011001100110011001100,
64'b0000111100001111111100001111000001101001100101100110100110010110,
64'b1100110000110011001100111100110010101010101010101010101010101010,
64'b0000111100001111111100001111000010101010010101010101010110101010,
64'b1100001100111100110000110011110000110011001100111100110011001100,
64'b0000000000000000000000000000000011001100110011001100110011001100,
64'b1100110011001100110011001100110001100110100110011001100101100110,
64'b1001100110011001011001100110011000111100110000111100001100111100,
64'b0011001100110011110011001100110010100101010110101010010101011010,
64'b0011001100110011110011001100110011111111000000001111111100000000,
64'b0101101010100101101001010101101011000011110000110011110000111100,
64'b0011110000111100001111000011110000001111111100000000111111110000,
64'b0011110000111100001111000011110000000000111111111111111100000000,
64'b0110011001100110011001100110011011110000111100001111000011110000,
64'b1111000011110000111100001111000010010110011010010110100110010110,
64'b0110011001100110011001100110011011001100110011001100110011001100,
64'b1100110000110011001100111100110000110011001100111100110011001100,
64'b0000000011111111111111110000000001011010010110100101101001011010,
64'b0000000000000000000000000000000001011010010110100101101001011010,
64'b1100110000110011001100111100110011000011110000110011110000111100,
64'b1111111100000000111111110000000001011010101001011010010101011010,
64'b1001100101100110100110010110011001100110100110011001100101100110,
64'b1001100101100110100110010110011011111111111111110000000000000000,
64'b1111111111111111000000000000000000001111111100000000111111110000,
64'b0110100110010110011010011001011010101010010101010101010110101010,
64'b1100001100111100110000110011110011111111111111110000000000000000,
64'b1001011010010110100101101001011001010101101010100101010110101010,
64'b1111111100000000111111110000000000111100110000111100001100111100,
64'b0011110000111100001111000011110001011010010110100101101001011010,
64'b0000111100001111111100001111000011110000111100001111000011110000,
64'b0101010101010101101010101010101010011001011001101001100101100110,
64'b1010101010101010101010101010101000110011110011000011001111001100,
64'b0000111100001111111100001111000000001111111100000000111111110000,
64'b0101010101010101101010101010101001100110100110011001100101100110,
64'b1100001111000011001111000011110001101001011010011001011010010110,
64'b1100001111000011001111000011110010101010101010101010101010101010,
64'b0000000000000000000000000000000010101010010101010101010110101010,
64'b1001011001101001011010011001011000110011001100111100110011001100,
64'b1111000000001111000011111111000010101010101010101010101010101010,
64'b1100001100111100110000110011110001100110011001100110011001100110,
64'b1111000000001111000011111111000001011010101001011010010101011010,
64'b1100110000110011001100111100110010011001011001101001100101100110,
64'b0110011010011001100110010110011011111111000000001111111100000000,
64'b0011110000111100001111000011110011000011110000110011110000111100,
64'b0110011001100110011001100110011000001111000011111111000011110000,
64'b1100001111000011001111000011110000000000111111111111111100000000,
64'b1010010101011010101001010101101011000011110000110011110000111100,
64'b0110011001100110011001100110011001101001100101100110100110010110,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b0011001111001100001100111100110000110011001100111100110011001100,
64'b1111000000001111000011111111000001011010010110100101101001011010,
64'b0110011010011001100110010110011001100110011001100110011001100110,
64'b0000111111110000000011111111000000111100001111000011110000111100,
64'b1010010110100101010110100101101011001100001100110011001111001100,
64'b0110011001100110011001100110011001101001011010011001011010010110,
64'b1111000011110000111100001111000011111111111111110000000000000000,
64'b1111111100000000111111110000000000001111111100000000111111110000,
64'b0011110000111100001111000011110001010101101010100101010110101010,
64'b0011001100110011110011001100110001010101010101011010101010101010,
64'b1010010110100101010110100101101010100101010110101010010101011010,
64'b1111111100000000111111110000000010010110011010010110100110010110,
64'b1111111100000000111111110000000000111100001111000011110000111100,
64'b1001011001101001011010011001011011110000111100001111000011110000,
64'b1100110000110011001100111100110010011001011001101001100101100110,
64'b1010010110100101010110100101101000111100001111000011110000111100,
64'b1111111100000000111111110000000000001111111100000000111111110000,
64'b1001100101100110100110010110011010101010010101010101010110101010,
64'b1001011010010110100101101001011010101010010101010101010110101010,
64'b1111111100000000111111110000000000110011001100111100110011001100,
64'b1111111111111111000000000000000011110000000011110000111111110000,
64'b0000111111110000000011111111000000110011001100111100110011001100,
64'b1111000011110000111100001111000011110000000011110000111111110000,
64'b1001100101100110100110010110011010100101101001010101101001011010,
64'b0101010101010101101010101010101011111111111111110000000000000000,
64'b1111111111111111000000000000000001100110011001100110011001100110,
64'b0011110011000011110000110011110001100110011001100110011001100110,
64'b1010010110100101010110100101101000001111000011111111000011110000,
64'b1001100101100110100110010110011011000011001111001100001100111100,
64'b1010101010101010101010101010101001010101101010100101010110101010,
64'b0110011010011001100110010110011000111100110000111100001100111100,
64'b0000000011111111111111110000000001011010010110100101101001011010,
64'b0110011001100110011001100110011011000011110000110011110000111100,
64'b0101101001011010010110100101101011110000000011110000111111110000,
64'b1010101001010101010101011010101001011010010110100101101001011010,
64'b1100001111000011001111000011110010010110100101101001011010010110,
64'b0000000011111111111111110000000001011010010110100101101001011010,
64'b0000111111110000000011111111000001101001100101100110100110010110,
64'b0110100110010110011010011001011001010101101010100101010110101010,
64'b1100001111000011001111000011110010100101010110101010010101011010,
64'b0101010110101010010101011010101000110011110011000011001111001100,
64'b1010010110100101010110100101101010010110011010010110100110010110,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b1100110000110011001100111100110001011010101001011010010101011010,
64'b1001011010010110100101101001011010011001011001101001100101100110,
64'b0000111100001111111100001111000000001111111100000000111111110000,
64'b0110100110010110011010011001011010101010010101010101010110101010,
64'b0011001100110011110011001100110010011001011001101001100101100110,
64'b1001100110011001011001100110011011000011001111001100001100111100,
64'b1001011001101001011010011001011000110011110011000011001111001100,
64'b0110100101101001100101101001011000111100110000111100001100111100,
64'b1111111111111111000000000000000000110011001100111100110011001100,
64'b1001011010010110100101101001011011001100001100110011001111001100,
64'b0101010101010101101010101010101000001111000011111111000011110000,
64'b1111111100000000111111110000000000111100110000111100001100111100,
64'b0011110000111100001111000011110010010110100101101001011010010110,
64'b1010010110100101010110100101101001100110100110011001100101100110,
64'b0110100110010110011010011001011001101001011010011001011010010110,
64'b1111111100000000111111110000000000000000111111111111111100000000,
64'b1001011001101001011010011001011000110011001100111100110011001100,
64'b1111000011110000111100001111000001101001011010011001011010010110,
64'b1001011010010110100101101001011011110000000011110000111111110000,
64'b1001011001101001011010011001011000001111000011111111000011110000,
64'b0110100110010110011010011001011011110000000011110000111111110000,
64'b1010101010101010101010101010101001011010010110100101101001011010,
64'b0110100110010110011010011001011010100101101001010101101001011010,
64'b1100110011001100110011001100110001010101101010100101010110101010,
64'b0101010101010101101010101010101001011010101001011010010101011010,
64'b0000111111110000000011111111000001101001100101100110100110010110,
64'b0011110000111100001111000011110001100110100110011001100101100110,
64'b0101010110101010010101011010101010101010010101010101010110101010,
64'b0110011001100110011001100110011011001100110011001100110011001100,
64'b0110011010011001100110010110011000000000000000000000000000000000,
64'b0101010110101010010101011010101001101001100101100110100110010110,
64'b1111111111111111000000000000000010010110100101101001011010010110,
64'b1111111111111111000000000000000010010110100101101001011010010110,
64'b0101010101010101101010101010101001101001011010011001011010010110,
64'b0000111111110000000011111111000001011010010110100101101001011010,
64'b1010010110100101010110100101101010101010101010101010101010101010,
64'b0011110000111100001111000011110001010101010101011010101010101010,
64'b0000000000000000000000000000000000000000111111111111111100000000,
64'b1111111100000000111111110000000011000011001111001100001100111100,
64'b0000000000000000000000000000000011000011110000110011110000111100,
64'b1111000011110000111100001111000010011001100110010110011001100110,
64'b1010010110100101010110100101101001011010010110100101101001011010,
64'b1001100110011001011001100110011000000000000000000000000000000000,
64'b1001100110011001011001100110011000111100110000111100001100111100,
64'b0011110011000011110000110011110011000011001111001100001100111100,
64'b0110100110010110011010011001011011000011001111001100001100111100,
64'b1010010101011010101001010101101011000011001111001100001100111100,
64'b0110100101101001100101101001011010011001011001101001100101100110,
64'b1010101010101010101010101010101011001100110011001100110011001100,
64'b0110100110010110011010011001011011001100110011001100110011001100,
64'b1100110011001100110011001100110001010101010101011010101010101010,
64'b1010101010101010101010101010101010100101010110101010010101011010,
64'b1010010101011010101001010101101000001111111100000000111111110000,
64'b0011110011000011110000110011110010010110100101101001011010010110,
64'b1010101001010101010101011010101010011001011001101001100101100110,
64'b1100110011001100110011001100110000000000000000000000000000000000,
64'b1001011010010110100101101001011011110000000011110000111111110000,
64'b0110011001100110011001100110011001011010101001011010010101011010,
64'b0101010101010101101010101010101011110000000011110000111111110000,
64'b0000111100001111111100001111000011110000000011110000111111110000,
64'b0000000000000000000000000000000011000011110000110011110000111100,
64'b1111111100000000111111110000000011110000111100001111000011110000,
64'b1111000000001111000011111111000011110000111100001111000011110000,
64'b0011110000111100001111000011110011001100110011001100110011001100,
64'b0110011001100110011001100110011010011001011001101001100101100110,
64'b0110011010011001100110010110011010101010010101010101010110101010,
64'b1111000000001111000011111111000011000011001111001100001100111100,
64'b1001100110011001011001100110011011000011110000110011110000111100,
64'b0101101001011010010110100101101000000000000000000000000000000000,
64'b1100001100111100110000110011110000000000111111111111111100000000,
64'b0011110000111100001111000011110001100110100110011001100101100110,
64'b1100110011001100110011001100110010101010010101010101010110101010,
64'b0101010110101010010101011010101010101010010101010101010110101010,
64'b1010101010101010101010101010101010100101010110101010010101011010,
64'b1111111111111111000000000000000001010101101010100101010110101010,
64'b0000000011111111111111110000000011111111000000001111111100000000,
64'b1010010101011010101001010101101011110000111100001111000011110000,
64'b0011110000111100001111000011110000111100001111000011110000111100,
64'b1100001111000011001111000011110010011001100110010110011001100110,
64'b1010101001010101010101011010101001011010101001011010010101011010,
64'b1001011010010110100101101001011000001111111100000000111111110000,
64'b1001100101100110100110010110011010101010101010101010101010101010,
64'b1111000000001111000011111111000011111111111111110000000000000000,
64'b0000111111110000000011111111000001101001011010011001011010010110,
64'b1111000011110000111100001111000010011001100110010110011001100110,
64'b0011001100110011110011001100110010011001100110010110011001100110,
64'b1100110011001100110011001100110001100110100110011001100101100110,
64'b0000000000000000000000000000000000110011001100111100110011001100,
64'b0101010101010101101010101010101011111111111111110000000000000000,
64'b0110011010011001100110010110011011111111000000001111111100000000,
64'b0000111111110000000011111111000000001111111100000000111111110000,
64'b1010010101011010101001010101101000111100001111000011110000111100,
64'b1001100110011001011001100110011001100110100110011001100101100110,
64'b0110100110010110011010011001011010101010010101010101010110101010,
64'b1100001111000011001111000011110011001100110011001100110011001100,
64'b0000000011111111111111110000000000000000000000000000000000000000,
64'b1010101001010101010101011010101001101001100101100110100110010110,
64'b1111111100000000111111110000000010010110100101101001011010010110,
64'b1111000011110000111100001111000010010110100101101001011010010110,
64'b0101101001011010010110100101101001101001011010011001011010010110,
64'b0000000000000000000000000000000001011010010110100101101001011010,
64'b1100110011001100110011001100110010101010101010101010101010101010,
64'b0110100101101001100101101001011001010101010101011010101010101010,
64'b0101010110101010010101011010101011111111000000001111111100000000,
64'b0110011010011001100110010110011011111111000000001111111100000000,
64'b1010010110100101010110100101101011000011001111001100001100111100,
64'b1111000011110000111100001111000011000011001111001100001100111100,
64'b0011110000111100001111000011110000110011110011000011001111001100,
64'b1100001111000011001111000011110001100110011001100110011001100110,
64'b1010010110100101010110100101101001011010101001011010010101011010,
64'b0011001100110011110011001100110010100101010110101010010101011010,
64'b1111000000001111000011111111000010101010101010101010101010101010,
64'b0000000011111111111111110000000001011010010110100101101001011010,
64'b0000000011111111111111110000000010101010101010101010101010101010,
64'b1001011010010110100101101001011010101010101010101010101010101010,
64'b1010101010101010101010101010101001101001100101100110100110010110,
64'b1111000011110000111100001111000011111111000000001111111100000000,
64'b1010010101011010101001010101101011111111111111110000000000000000,
64'b0011110011000011110000110011110011110000000011110000111111110000,
64'b1010010101011010101001010101101011110000000011110000111111110000,
64'b0011001111001100001100111100110000001111000011111111000011110000,
64'b1100110000110011001100111100110000111100001111000011110000111100,
64'b0011110011000011110000110011110011001100001100110011001111001100,
64'b0110100101101001100101101001011001100110100110011001100101100110,
64'b0101101001011010010110100101101011001100110011001100110011001100,
64'b0101010110101010010101011010101000110011110011000011001111001100,
64'b0101010110101010010101011010101011001100110011001100110011001100,
64'b1111111100000000111111110000000011001100110011001100110011001100,
64'b0110011001100110011001100110011000111100110000111100001100111100,
64'b0000111111110000000011111111000000000000000000000000000000000000,
64'b1010101010101010101010101010101000000000000000000000000000000000,
64'b0101010110101010010101011010101010101010010101010101010110101010,
64'b1001011001101001011010011001011010101010010101010101010110101010,
64'b0011001100110011110011001100110001010101101010100101010110101010,
64'b1100110011001100110011001100110010100101010110101010010101011010,
64'b1111111100000000111111110000000000001111000011111111000011110000,
64'b0101101010100101101001010101101001101001011010011001011010010110,
64'b0110100101101001100101101001011001011010010110100101101001011010,
64'b0011001111001100001100111100110000001111000011111111000011110000,
64'b0011001111001100001100111100110011110000111100001111000011110000,
64'b0110100101101001100101101001011011110000111100001111000011110000,
64'b1001011010010110100101101001011011110000000011110000111111110000,
64'b0000111111110000000011111111000010101010101010101010101010101010,
64'b1100110011001100110011001100110010101010101010101010101010101010,
64'b0011001100110011110011001100110000110011001100111100110011001100,
64'b0011110011000011110000110011110010011001100110010110011001100110,
64'b0101101001011010010110100101101010011001100110010110011001100110,
64'b0101101001011010010110100101101011001100001100110011001111001100,
64'b1111111111111111000000000000000011111111000000001111111100000000,
64'b1100110000110011001100111100110001101001100101100110100110010110,
64'b0110100110010110011010011001011010011001011001101001100101100110,
64'b1010010110100101010110100101101011111111000000001111111100000000,
64'b0000111100001111111100001111000001010101101010100101010110101010,
64'b1100001100111100110000110011110011111111000000001111111100000000,
64'b0110100110010110011010011001011000000000111111111111111100000000,
64'b1111111100000000111111110000000001100110011001100110011001100110,
64'b0011110011000011110000110011110011001100110011001100110011001100,
64'b0101010101010101101010101010101011110000111100001111000011110000,
64'b1010101001010101010101011010101010010110100101101001011010010110,
64'b1010010101011010101001010101101010010110100101101001011010010110,
64'b1111000000001111000011111111000010100101101001010101101001011010,
64'b1010010110100101010110100101101001010101010101011010101010101010,
64'b1001011010010110100101101001011000111100110000111100001100111100,
64'b0110011001100110011001100110011011000011110000110011110000111100,
64'b0011001100110011110011001100110011111111111111110000000000000000,
64'b0101010101010101101010101010101000110011001100111100110011001100,
64'b1100110000110011001100111100110011111111111111110000000000000000,
64'b1001011001101001011010011001011011111111111111110000000000000000,
64'b1111000011110000111100001111000010010110100101101001011010010110,
64'b0011110000111100001111000011110011110000111100001111000011110000,
64'b1100001111000011001111000011110011111111000000001111111100000000,
64'b0110100101101001100101101001011011000011001111001100001100111100,
64'b0101101010100101101001010101101011000011001111001100001100111100,
64'b1100001100111100110000110011110000110011110011000011001111001100,
64'b0011110011000011110000110011110001100110011001100110011001100110,
64'b0101101010100101101001010101101001011010101001011010010101011010,
64'b1100110000110011001100111100110010100101010110101010010101011010,
64'b1111000000001111000011111111000010101010101010101010101010101010,
64'b0110011010011001100110010110011001011010010110100101101001011010,
64'b0011001100110011110011001100110010101010101010101010101010101010,
64'b0011110011000011110000110011110010101010101010101010101010101010,
64'b1010010101011010101001010101101001101001100101100110100110010110,
64'b1010010101011010101001010101101000110011001100111100110011001100,
64'b0000111111110000000011111111000001011010010110100101101001011010,
64'b0110100110010110011010011001011000000000111111111111111100000000,
64'b0110011010011001100110010110011011001100001100110011001111001100,
64'b0101101010100101101001010101101011001100110011001100110011001100,
64'b1111000000001111000011111111000010011001100110010110011001100110,
64'b0110011010011001100110010110011011111111000000001111111100000000,
64'b1010010110100101010110100101101010010110100101101001011010010110,
64'b1010101001010101010101011010101011001100001100110011001111001100,
64'b0110100101101001100101101001011000110011001100111100110011001100,
64'b0101101001011010010110100101101001011010010110100101101001011010,
64'b0101101010100101101001010101101001100110011001100110011001100110,
64'b1001100101100110100110010110011000110011110011000011001111001100,
64'b1010101010101010101010101010101000111100110000111100001100111100,
64'b1010010101011010101001010101101000111100110000111100001100111100,
64'b1100110000110011001100111100110000001111000011111111000011110000,
64'b1111111111111111000000000000000010011001100110010110011001100110,
64'b1010010101011010101001010101101010011001100110010110011001100110,
64'b0000111111110000000011111111000010011001100110010110011001100110,
64'b0101101001011010010110100101101001100110011001100110011001100110,
64'b0110100101101001100101101001011000110011001100111100110011001100,
64'b1001100101100110100110010110011000001111111100000000111111110000,
64'b0110100101101001100101101001011001011010101001011010010101011010,
64'b0000111111110000000011111111000000001111111100000000111111110000,
64'b0110011010011001100110010110011010010110100101101001011010010110,
64'b0110011001100110011001100110011000000000000000000000000000000000,
64'b1010101001010101010101011010101011110000000011110000111111110000,
64'b0110100110010110011010011001011001011010101001011010010101011010,
64'b1111111111111111000000000000000001010101101010100101010110101010,
64'b1001011010010110100101101001011010010110100101101001011010010110,
64'b1010010101011010101001010101101010010110100101101001011010010110,
64'b1010010101011010101001010101101010010110100101101001011010010110,
64'b0000000011111111111111110000000010010110100101101001011010010110,
64'b0011001100110011110011001100110011110000111100001111000011110000,
64'b0110100110010110011010011001011010101010010101010101010110101010,
64'b1100001111000011001111000011110011001100001100110011001111001100,
64'b0011110011000011110000110011110010101010010101010101010110101010,
64'b0110100101101001100101101001011011000011001111001100001100111100,
64'b0110011001100110011001100110011000000000000000000000000000000000,
64'b0011001100110011110011001100110000000000111111111111111100000000,
64'b1001011001101001011010011001011001100110100110011001100101100110,
64'b0000000000000000000000000000000010011001100110010110011001100110,
64'b0110100110010110011010011001011011000011001111001100001100111100,
64'b1100110000110011001100111100110011000011001111001100001100111100,
64'b1100110000110011001100111100110011000011001111001100001100111100,
64'b1111111111111111000000000000000011000011001111001100001100111100,
64'b0101101001011010010110100101101011111111000000001111111100000000,
64'b1001011001101001011010011001011000110011001100111100110011001100,
64'b0000111111110000000011111111000010100101101001010101101001011010,
64'b0101101010100101101001010101101010011001100110010110011001100110,
64'b0110100110010110011010011001011001011010101001011010010101011010,
64'b1001011010010110100101101001011000000000000000000000000000000000,
64'b0011110011000011110000110011110000110011110011000011001111001100,
64'b0011001111001100001100111100110011001100110011001100110011001100,
64'b0101101001011010010110100101101001100110011001100110011001100110,
64'b0000000011111111111111110000000001100110100110011001100101100110,
64'b1100110011001100110011001100110000110011110011000011001111001100,
64'b0000000000000000000000000000000001010101101010100101010110101010,
64'b1001100110011001011001100110011011000011001111001100001100111100,
64'b0110100101101001100101101001011000001111111100000000111111110000,
64'b0011110000111100001111000011110011110000000011110000111111110000,
64'b1010101010101010101010101010101010011001100110010110011001100110,
64'b0101101010100101101001010101101000000000000000000000000000000000,
64'b0011110011000011110000110011110011001100001100110011001111001100,
64'b0011001111001100001100111100110001011010010110100101101001011010,
64'b0011110000111100001111000011110010100101101001010101101001011010,
64'b0000000000000000000000000000000011110000111100001111000011110000,
64'b1100001100111100110000110011110000111100001111000011110000111100,
64'b1100001111000011001111000011110011000011110000110011110000111100,
64'b1001100110011001011001100110011010100101101001010101101001011010,
64'b1010010110100101010110100101101000110011001100111100110011001100,
64'b0000111100001111111100001111000011110000000011110000111111110000,
64'b1001100110011001011001100110011000000000111111111111111100000000,
64'b1010010110100101010110100101101000000000111111111111111100000000,
64'b1100110000110011001100111100110010010110100101101001011010010110,
64'b0101101010100101101001010101101010101010101010101010101010101010,
64'b1111000000001111000011111111000000001111000011111111000011110000,
64'b1010101010101010101010101010101010011001011001101001100101100110,
64'b0110100101101001100101101001011010011001011001101001100101100110,
64'b1010010110100101010110100101101001010101101010100101010110101010,
64'b0000000011111111111111110000000000001111111100000000111111110000,
64'b0011001111001100001100111100110000001111111100000000111111110000,
64'b0101010101010101101010101010101010011001011001101001100101100110,
64'b0011110011000011110000110011110001011010010110100101101001011010,
64'b0110011010011001100110010110011010101010010101010101010110101010,
64'b0110011010011001100110010110011001010101010101011010101010101010,
64'b1001100110011001011001100110011001010101010101011010101010101010,
64'b1010010101011010101001010101101001101001100101100110100110010110,
64'b1111000000001111000011111111000011001100110011001100110011001100,
64'b0000000011111111111111110000000011111111000000001111111100000000,
64'b1001011010010110100101101001011010010110100101101001011010010110,
64'b1100001100111100110000110011110001101001011010011001011010010110,
64'b1001100101100110100110010110011000110011001100111100110011001100,
64'b0101010101010101101010101010101000000000111111111111111100000000,
64'b1010010110100101010110100101101000000000111111111111111100000000,
64'b1100110011001100110011001100110011000011110000110011110000111100,
64'b0101101010100101101001010101101000110011110011000011001111001100,
64'b0110100101101001100101101001011000110011001100111100110011001100,
64'b0110100101101001100101101001011001100110011001100110011001100110,
64'b1001011010010110100101101001011001100110011001100110011001100110,
64'b0110011010011001100110010110011010010110011010010110100110010110,
64'b0000000011111111111111110000000011110000111100001111000011110000,
64'b0101010101010101101010101010101011111111111111110000000000000000,
64'b0110100110010110011010011001011011000011001111001100001100111100,
64'b1111000000001111000011111111000011000011001111001100001100111100,
64'b1100001111000011001111000011110001011010010110100101101001011010,
64'b1100110011001100110011001100110001010101010101011010101010101010,
64'b1001100101100110100110010110011001010101010101011010101010101010,
64'b0101101001011010010110100101101010100101010110101010010101011010,
64'b1100110000110011001100111100110010100101101001010101101001011010,
64'b0110100110010110011010011001011011110000111100001111000011110000,
64'b0110100110010110011010011001011010010110100101101001011010010110,
64'b0110100110010110011010011001011000111100001111000011110000111100,
64'b1100001111000011001111000011110000111100110000111100001100111100,
64'b0101010101010101101010101010101001010101101010100101010110101010,
64'b0110011001100110011001100110011000000000000000000000000000000000,
64'b0110100110010110011010011001011010100101010110101010010101011010,
64'b1010101001010101010101011010101001011010101001011010010101011010,
64'b1010010101011010101001010101101000110011110011000011001111001100,
64'b0101101001011010010110100101101011001100110011001100110011001100,
64'b1100001111000011001111000011110001100110011001100110011001100110,
64'b0011001111001100001100111100110001100110100110011001100101100110,
64'b0000111100001111111100001111000000110011110011000011001111001100,
64'b1001011001101001011010011001011001010101101010100101010110101010,
64'b0011110011000011110000110011110011000011001111001100001100111100,
64'b0011110011000011110000110011110000001111111100000000111111110000,
64'b0000111111110000000011111111000011110000000011110000111111110000,
64'b0110011001100110011001100110011010011001100110010110011001100110,
64'b1001011010010110100101101001011000000000000000000000000000000000,
64'b1100001100111100110000110011110000110011110011000011001111001100,
64'b0110100101101001100101101001011000000000000000000000000000000000,
64'b1100001100111100110000110011110001011010010110100101101001011010,
64'b0000000000000000000000000000000010100101101001010101101001011010,
64'b1111111100000000111111110000000010101010010101010101010110101010,
64'b1100110000110011001100111100110010011001100110010110011001100110,
64'b0011001100110011110011001100110001101001011010011001011010010110,
64'b1010101010101010101010101010101010100101101001010101101001011010,
64'b0110100110010110011010011001011001011010010110100101101001011010,
64'b0000000000000000000000000000000010100101101001010101101001011010,
64'b0110011001100110011001100110011010010110100101101001011010010110,
64'b0101101010100101101001010101101011000011110000110011110000111100,
64'b1100110011001100110011001100110011111111000000001111111100000000,
64'b0101010110101010010101011010101000001111111100000000111111110000,
64'b1010101001010101010101011010101010101010101010101010101010101010,
64'b1001100110011001011001100110011000110011110011000011001111001100,
64'b0000000000000000000000000000000000110011110011000011001111001100,
64'b0000000011111111111111110000000010011001100110010110011001100110,
64'b1100001100111100110000110011110010010110100101101001011010010110,
64'b0110100101101001100101101001011001101001100101100110100110010110,
64'b1100110011001100110011001100110010011001011001101001100101100110,
64'b0101010101010101101010101010101010011001011001101001100101100110,
64'b0000000000000000000000000000000000110011110011000011001111001100,
64'b0101101001011010010110100101101001101001100101100110100110010110,
64'b1001011010010110100101101001011000001111111100000000111111110000,
64'b1001011010010110100101101001011001010101010101011010101010101010,
64'b1001100101100110100110010110011011111111000000001111111100000000,
64'b1111000011110000111100001111000011001100110011001100110011001100,
64'b0101010110101010010101011010101000001111000011111111000011110000,
64'b1010101010101010101010101010101000001111000011111111000011110000,
64'b0000000011111111111111110000000000111100001111000011110000111100,
64'b1001011010010110100101101001011001101001100101100110100110010110,
64'b1111000000001111000011111111000000111100110000111100001100111100,
64'b1111000011110000111100001111000011000011110000110011110000111100,
64'b1010010101011010101001010101101011000011110000110011110000111100,
64'b1010101010101010101010101010101000001111000011111111000011110000,
64'b0101010110101010010101011010101000111100110000111100001100111100,
64'b1001100110011001011001100110011000000000111111111111111100000000,
64'b0000111111110000000011111111000011001100110011001100110011001100,
64'b0110100110010110011010011001011010101010101010101010101010101010,
64'b0101010110101010010101011010101011110000111100001111000011110000,
64'b0011001100110011110011001100110011111111000000001111111100000000,
64'b1100110011001100110011001100110001010101101010100101010110101010,
64'b1111111111111111000000000000000010100101010110101010010101011010,
64'b0110100110010110011010011001011000111100110000111100001100111100,
64'b0000000011111111111111110000000011110000000011110000111111110000,
64'b0101010110101010010101011010101010100101010110101010010101011010,
64'b1100110000110011001100111100110010100101010110101010010101011010,
64'b1100110011001100110011001100110001010101101010100101010110101010,
64'b0011001100110011110011001100110001011010101001011010010101011010,
64'b0011110000111100001111000011110001010101010101011010101010101010,
64'b1010101001010101010101011010101001011010010110100101101001011010,
64'b1100001100111100110000110011110011001100110011001100110011001100,
64'b1111000011110000111100001111000011111111000000001111111100000000,
64'b0011001111001100001100111100110011111111111111110000000000000000,
64'b0101101001011010010110100101101000110011001100111100110011001100,
64'b1111111100000000111111110000000011001100001100110011001111001100,
64'b0101101001011010010110100101101011110000000011110000111111110000,
64'b1100110011001100110011001100110010101010010101010101010110101010,
64'b0011001100110011110011001100110001100110100110011001100101100110,
64'b0110011010011001100110010110011011001100001100110011001111001100,
64'b0101101001011010010110100101101000110011001100111100110011001100,
64'b1001011010010110100101101001011011001100001100110011001111001100,
64'b1111111111111111000000000000000001100110011001100110011001100110,
64'b1111111111111111000000000000000010011001011001101001100101100110,
64'b1111000011110000111100001111000011110000111100001111000011110000,
64'b1001011001101001011010011001011011111111111111110000000000000000,
64'b1100110000110011001100111100110000000000000000000000000000000000,
64'b0011001111001100001100111100110001011010010110100101101001011010,
64'b0000000011111111111111110000000010100101101001010101101001011010,
64'b1111111111111111000000000000000010101010010101010101010110101010,
64'b1100001111000011001111000011110010011001100110010110011001100110,
64'b0101101001011010010110100101101001101001011010011001011010010110,
64'b0000000011111111111111110000000010100101101001010101101001011010,
64'b1001100101100110100110010110011001011010010110100101101001011010,
64'b1010010101011010101001010101101010100101101001010101101001011010,
64'b0101101010100101101001010101101010010110100101101001011010010110,
64'b0110011001100110011001100110011011000011110000110011110000111100,
64'b0000000000000000000000000000000011111111000000001111111100000000,
64'b1001011001101001011010011001011011000011110000110011110000111100,
64'b1010010110100101010110100101101001101001100101100110100110010110,
64'b1010010110100101010110100101101000110011110011000011001111001100,
64'b1111111111111111000000000000000011001100110011001100110011001100,
64'b1010101010101010101010101010101001010101101010100101010110101010,
64'b1010010101011010101001010101101010100101101001010101101001011010,
64'b1001100101100110100110010110011011000011001111001100001100111100,
64'b1111111111111111000000000000000011110000111100001111000011110000,
64'b0110100101101001100101101001011010011001011001101001100101100110,
64'b1100110000110011001100111100110001010101101010100101010110101010,
64'b1100110000110011001100111100110000110011001100111100110011001100,
64'b1001011010010110100101101001011011000011001111001100001100111100,
64'b0000000000000000000000000000000011111111000000001111111100000000,
64'b1111111100000000111111110000000011001100001100110011001111001100,
64'b0101101001011010010110100101101001010101010101011010101010101010,
64'b1001100101100110100110010110011000001111000011111111000011110000,
64'b0101010110101010010101011010101000001111111100000000111111110000,
64'b1010101001010101010101011010101011111111000000001111111100000000,
64'b1111111100000000111111110000000000000000111111111111111100000000,
64'b0110100101101001100101101001011011110000000011110000111111110000,
64'b0110100110010110011010011001011010010110100101101001011010010110,
64'b0110100110010110011010011001011011000011110000110011110000111100,
64'b1100001111000011001111000011110001010101010101011010101010101010,
64'b1111111100000000111111110000000010101010010101010101010110101010,
64'b1010010101011010101001010101101010010110011010010110100110010110,
64'b0101010110101010010101011010101001010101101010100101010110101010,
64'b1001011010010110100101101001011000001111000011111111000011110000,
64'b1111000011110000111100001111000001100110011001100110011001100110,
64'b1100001111000011001111000011110001010101101010100101010110101010,
64'b1100110000110011001100111100110010101010010101010101010110101010,
64'b1111111100000000111111110000000011111111111111110000000000000000,
64'b0110011001100110011001100110011011111111111111110000000000000000,
64'b0110100110010110011010011001011010101010010101010101010110101010,
64'b1111111111111111000000000000000001101001100101100110100110010110,
64'b0011110011000011110000110011110000001111111100000000111111110000,
64'b0110100110010110011010011001011001100110011001100110011001100110,
64'b0000111111110000000011111111000010011001100110010110011001100110,
64'b0000000011111111111111110000000010010110011010010110100110010110,
64'b1001100101100110100110010110011001100110011001100110011001100110,
64'b1100001100111100110000110011110011111111000000001111111100000000,
64'b1111111100000000111111110000000010010110100101101001011010010110,
64'b0000111111110000000011111111000000110011001100111100110011001100,
64'b1010010110100101010110100101101000110011001100111100110011001100,
64'b0101010101010101101010101010101010101010101010101010101010101010,
64'b0011110000111100001111000011110010101010101010101010101010101010,
64'b0011110011000011110000110011110010011001100110010110011001100110,
64'b0000000000000000000000000000000010010110011010010110100110010110,
64'b0101101010100101101001010101101000000000111111111111111100000000,
64'b1001011001101001011010011001011000111100001111000011110000111100,
64'b0000000011111111111111110000000000111100001111000011110000111100,
64'b1111111111111111000000000000000010010110011010010110100110010110,
64'b1001011010010110100101101001011010010110100101101001011010010110,
64'b1001100101100110100110010110011010010110100101101001011010010110,
64'b0011110011000011110000110011110000000000000000000000000000000000,
64'b0000000011111111111111110000000011110000111100001111000011110000,
64'b1100110011001100110011001100110010100101010110101010010101011010,
64'b1010101001010101010101011010101010101010010101010101010110101010,
64'b1001011001101001011010011001011011111111111111110000000000000000,
64'b0101101010100101101001010101101010010110100101101001011010010110,
64'b1100001100111100110000110011110011111111111111110000000000000000,
64'b1100110000110011001100111100110001010101010101011010101010101010,
64'b1111000000001111000011111111000011000011001111001100001100111100,
64'b0000111111110000000011111111000001010101010101011010101010101010,
64'b0110011001100110011001100110011011110000000011110000111111110000,
64'b0011110000111100001111000011110000111100001111000011110000111100,
64'b0000000000000000000000000000000011000011001111001100001100111100,
64'b0011001100110011110011001100110000000000000000000000000000000000,
64'b0101010101010101101010101010101011111111000000001111111100000000,
64'b1010010101011010101001010101101011001100001100110011001111001100,
64'b1111111100000000111111110000000000110011001100111100110011001100,
64'b1010010101011010101001010101101010101010101010101010101010101010,
64'b1100110000110011001100111100110001101001100101100110100110010110,
64'b0011001100110011110011001100110000000000000000000000000000000000,
64'b0000111100001111111100001111000001100110011001100110011001100110,
64'b1100110000110011001100111100110001011010101001011010010101011010,
64'b1111000011110000111100001111000011001100110011001100110011001100,
64'b1111000011110000111100001111000010101010010101010101010110101010,
64'b0101101001011010010110100101101010100101010110101010010101011010,
64'b0110100101101001100101101001011001011010101001011010010101011010,
64'b0011001111001100001100111100110000000000000000000000000000000000,
64'b0110011001100110011001100110011011111111111111110000000000000000,
64'b1001100110011001011001100110011000001111000011111111000011110000,
64'b0011001111001100001100111100110001011010010110100101101001011010,
64'b1111111100000000111111110000000001100110011001100110011001100110,
64'b1010010110100101010110100101101000111100110000111100001100111100,
64'b0011001111001100001100111100110000000000000000000000000000000000,
64'b0101010110101010010101011010101000111100001111000011110000111100,
64'b1100001111000011001111000011110011001100001100110011001111001100,
64'b0000111100001111111100001111000001011010010110100101101001011010,
64'b0011001111001100001100111100110000110011001100111100110011001100,
64'b0110011001100110011001100110011010011001011001101001100101100110,
64'b1100001100111100110000110011110011001100001100110011001111001100,
64'b1010010110100101010110100101101010101010101010101010101010101010,
64'b0011110000111100001111000011110000000000000000000000000000000000,
64'b0011110000111100001111000011110001010101101010100101010110101010,
64'b1010010110100101010110100101101010011001011001101001100101100110,
64'b1111111111111111000000000000000000111100001111000011110000111100,
64'b0011001111001100001100111100110011110000000011110000111111110000,
64'b1010010110100101010110100101101010101010101010101010101010101010,
64'b0011001100110011110011001100110000001111111100000000111111110000,
64'b0000111111110000000011111111000000001111000011111111000011110000,
64'b0101010110101010010101011010101010011001011001101001100101100110,
64'b1010010110100101010110100101101011110000111100001111000011110000,
64'b0011110000111100001111000011110010010110100101101001011010010110,
64'b0101101010100101101001010101101010100101101001010101101001011010,
64'b0011001111001100001100111100110001100110011001100110011001100110,
64'b1010010101011010101001010101101000000000000000000000000000000000,
64'b0000111111110000000011111111000000110011001100111100110011001100,
64'b0011001111001100001100111100110011000011110000110011110000111100,
64'b1010101010101010101010101010101000001111111100000000111111110000,
64'b1010010110100101010110100101101000000000111111111111111100000000,
64'b0011001111001100001100111100110001100110011001100110011001100110,
64'b0101101001011010010110100101101000000000111111111111111100000000,
64'b1010101001010101010101011010101011111111000000001111111100000000,
64'b0011001100110011110011001100110001101001011010011001011010010110,
64'b0011001111001100001100111100110011111111000000001111111100000000,
64'b1010010101011010101001010101101011000011001111001100001100111100,
64'b0110011010011001100110010110011010011001011001101001100101100110,
64'b1010010110100101010110100101101010010110100101101001011010010110,
64'b1100110000110011001100111100110000000000000000000000000000000000,
64'b0000000011111111111111110000000011110000111100001111000011110000,
64'b0000111100001111111100001111000010100101010110101010010101011010,
64'b1100110011001100110011001100110010101010010101010101010110101010,
64'b0011001111001100001100111100110011111111111111110000000000000000,
64'b1010010110100101010110100101101010010110100101101001011010010110,
64'b0011001111001100001100111100110011111111111111110000000000000000,
64'b0011001100110011110011001100110001010101010101011010101010101010,
64'b0101101001011010010110100101101011000011001111001100001100111100,
64'b1010010110100101010110100101101001010101010101011010101010101010,
64'b0011001111001100001100111100110000001111111100000000111111110000,
64'b0110011010011001100110010110011011111111000000001111111100000000,
64'b0011110011000011110000110011110011001100001100110011001111001100,
64'b1100110000110011001100111100110001100110100110011001100101100110,
64'b1010010110100101010110100101101000000000111111111111111100000000,
64'b0000000011111111111111110000000010100101010110101010010101011010,
64'b1010101001010101010101011010101010100101010110101010010101011010,
64'b0011110000111100001111000011110010100101101001010101101001011010,
64'b0110011001100110011001100110011000000000000000000000000000000000,
64'b0101010110101010010101011010101010010110100101101001011010010110,
64'b0011001111001100001100111100110000111100110000111100001100111100,
64'b0000000011111111111111110000000001101001011010011001011010010110,
64'b0101010101010101101010101010101000000000000000000000000000000000,
64'b1001100101100110100110010110011001010101101010100101010110101010,
64'b0000111111110000000011111111000001010101010101011010101010101010,
64'b0110011001100110011001100110011000001111000011111111000011110000,
64'b0110100110010110011010011001011001101001011010011001011010010110,
64'b0011110011000011110000110011110001010101010101011010101010101010,
64'b0101010110101010010101011010101001100110100110011001100101100110,
64'b0011001111001100001100111100110011001100001100110011001111001100,
64'b1001100101100110100110010110011000110011110011000011001111001100,
64'b0101101001011010010110100101101010101010101010101010101010101010,
64'b0110011010011001100110010110011011000011001111001100001100111100,
64'b0011110011000011110000110011110011110000000011110000111111110000,
64'b1111111100000000111111110000000001101001100101100110100110010110,
64'b0011001100110011110011001100110010101010101010101010101010101010,
64'b0000111111110000000011111111000011001100110011001100110011001100,
64'b1100110011001100110011001100110001100110011001100110011001100110,
64'b0000000011111111111111110000000001010101101010100101010110101010,
64'b1111000011110000111100001111000001101001100101100110100110010110,
64'b0101010110101010010101011010101001100110011001100110011001100110,
64'b1001100101100110100110010110011001101001011010011001011010010110,
64'b1010010101011010101001010101101010100101101001010101101001011010,
64'b1111111111111111000000000000000010100101101001010101101001011010,
64'b0101010110101010010101011010101011001100110011001100110011001100,
64'b1001011001101001011010011001011011110000000011110000111111110000,
64'b0110100101101001100101101001011000000000111111111111111100000000,
64'b0101010110101010010101011010101010010110011010010110100110010110,
64'b1010010110100101010110100101101011001100110011001100110011001100,
64'b1100110011001100110011001100110011110000111100001111000011110000,
64'b0101101001011010010110100101101000111100001111000011110000111100,
64'b1111111111111111000000000000000000110011001100111100110011001100,
64'b0101010110101010010101011010101000111100110000111100001100111100,
64'b0011001100110011110011001100110000111100001111000011110000111100,
64'b1100001111000011001111000011110011000011001111001100001100111100,
64'b1100110000110011001100111100110010011001011001101001100101100110,
64'b0000000000000000000000000000000010011001011001101001100101100110,
64'b1001100110011001011001100110011001011010010110100101101001011010,
64'b0011110011000011110000110011110000000000111111111111111100000000,
64'b0110100110010110011010011001011001010101010101011010101010101010,
64'b1001100110011001011001100110011010010110011010010110100110010110,
64'b0011001111001100001100111100110001011010010110100101101001011010,
64'b0101101001011010010110100101101011111111000000001111111100000000,
64'b1111111111111111000000000000000000001111111100000000111111110000,
64'b0011110011000011110000110011110011110000111100001111000011110000,
64'b0101010110101010010101011010101001011010101001011010010101011010,
64'b0101010101010101101010101010101010100101010110101010010101011010,
64'b1010010110100101010110100101101011110000000011110000111111110000,
64'b0000111111110000000011111111000011000011110000110011110000111100,
64'b1001011010010110100101101001011011000011110000110011110000111100,
64'b0101101001011010010110100101101000110011110011000011001111001100,
64'b0000111100001111111100001111000011111111111111110000000000000000,
64'b1010010110100101010110100101101001100110011001100110011001100110,
64'b0011110011000011110000110011110010010110011010010110100110010110,
64'b1111000011110000111100001111000010011001011001101001100101100110,
64'b1010101010101010101010101010101000000000000000000000000000000000,
64'b0110011010011001100110010110011000000000111111111111111100000000,
64'b0110011001100110011001100110011011111111000000001111111100000000,
64'b0101010110101010010101011010101011001100001100110011001111001100,
64'b0110100101101001100101101001011001100110100110011001100101100110,
64'b1001100110011001011001100110011000000000111111111111111100000000,
64'b0000000000000000000000000000000010100101010110101010010101011010,
64'b1111111100000000111111110000000010100101010110101010010101011010,
64'b0101010110101010010101011010101010100101101001010101101001011010,
64'b1010101010101010101010101010101000000000000000000000000000000000,
64'b1010101010101010101010101010101010010110100101101001011010010110,
64'b0101101001011010010110100101101000111100110000111100001100111100,
64'b0000000011111111111111110000000001101001011010011001011010010110,
64'b0101010110101010010101011010101000000000000000000000000000000000,
64'b1100001111000011001111000011110000110011110011000011001111001100,
64'b1001011010010110100101101001011001101001100101100110100110010110,
64'b0011001100110011110011001100110011000011001111001100001100111100,
64'b1100001100111100110000110011110011001100110011001100110011001100,
64'b1001011010010110100101101001011001010101101010100101010110101010,
64'b1010101010101010101010101010101011001100110011001100110011001100,
64'b1111111111111111000000000000000011110000000011110000111111110000,
64'b0011001100110011110011001100110001010101101010100101010110101010,
64'b1100110011001100110011001100110011111111000000001111111100000000,
64'b1100110011001100110011001100110011110000111100001111000011110000,
64'b0011001111001100001100111100110011110000111100001111000011110000,
64'b1111111111111111000000000000000000111100110000111100001100111100,
64'b0110011001100110011001100110011000110011110011000011001111001100,
64'b0110100101101001100101101001011011000011001111001100001100111100,
64'b0101010101010101101010101010101000000000000000000000000000000000,
64'b0011110011000011110000110011110000111100001111000011110000111100,
64'b1111111100000000111111110000000001010101010101011010101010101010,
64'b1100001111000011001111000011110000110011110011000011001111001100,
64'b0110011010011001100110010110011001011010101001011010010101011010,
64'b0011110000111100001111000011110000111100110000111100001100111100,
64'b0011110000111100001111000011110011111111111111110000000000000000,
64'b0000111111110000000011111111000010101010010101010101010110101010,
64'b1100001100111100110000110011110011001100110011001100110011001100,
64'b0000111111110000000011111111000011111111111111110000000000000000,
64'b0101010101010101101010101010101010100101010110101010010101011010,
64'b0000111111110000000011111111000011000011001111001100001100111100,
64'b0000111100001111111100001111000001011010101001011010010101011010,
64'b0101101010100101101001010101101000000000000000000000000000000000,
64'b1001011010010110100101101001011000001111111100000000111111110000,
64'b1111000011110000111100001111000011001100110011001100110011001100,
64'b0000111100001111111100001111000010100101101001010101101001011010,
64'b1100001100111100110000110011110011001100001100110011001111001100,
64'b1001100101100110100110010110011001011010101001011010010101011010,
64'b0110100110010110011010011001011010101010101010101010101010101010,
64'b0101010101010101101010101010101010011001100110010110011001100110,
64'b1100001111000011001111000011110001011010010110100101101001011010,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1001100110011001011001100110011001100110100110011001100101100110,
64'b1100110011001100110011001100110000001111111100000000111111110000,
64'b0101010110101010010101011010101011001100001100110011001111001100,
64'b0110011010011001100110010110011010101010101010101010101010101010,
64'b0110100110010110011010011001011000000000111111111111111100000000,
64'b1111111100000000111111110000000011110000111100001111000011110000,
64'b1111111100000000111111110000000000110011110011000011001111001100,
64'b0101101010100101101001010101101010100101101001010101101001011010,
64'b1100001111000011001111000011110001100110100110011001100101100110,
64'b0011110011000011110000110011110001100110011001100110011001100110,
64'b1100110011001100110011001100110000111100001111000011110000111100,
64'b1010010101011010101001010101101010011001011001101001100101100110,
64'b1010101010101010101010101010101000000000000000000000000000000000,
64'b0011110000111100001111000011110011000011110000110011110000111100,
64'b0101101001011010010110100101101001010101101010100101010110101010,
64'b0101010110101010010101011010101001101001100101100110100110010110,
64'b1111111100000000111111110000000001011010101001011010010101011010,
64'b0101101001011010010110100101101000110011110011000011001111001100,
64'b0101101001011010010110100101101011110000000011110000111111110000,
64'b1111111100000000111111110000000000001111111100000000111111110000,
64'b0110011001100110011001100110011010011001100110010110011001100110,
64'b1001100101100110100110010110011001010101010101011010101010101010,
64'b0011110011000011110000110011110011110000111100001111000011110000,
64'b0000111111110000000011111111000001011010010110100101101001011010,
64'b1111111111111111000000000000000011110000000011110000111111110000,
64'b1100110000110011001100111100110000000000111111111111111100000000,
64'b0101101010100101101001010101101001011010101001011010010101011010,
64'b1010101010101010101010101010101011111111000000001111111100000000,
64'b0101010110101010010101011010101000111100110000111100001100111100,
64'b1100001100111100110000110011110011001100001100110011001111001100,
64'b1111111111111111000000000000000010100101101001010101101001011010,
64'b1001011001101001011010011001011000000000111111111111111100000000,
64'b1111111100000000111111110000000010101010010101010101010110101010,
64'b1001011001101001011010011001011000111100001111000011110000111100,
64'b1111111111111111000000000000000001100110011001100110011001100110,
64'b1001011001101001011010011001011001010101101010100101010110101010,
64'b1111111111111111000000000000000000110011110011000011001111001100,
64'b0011001111001100001100111100110000000000111111111111111100000000,
64'b1010010101011010101001010101101001010101010101011010101010101010,
64'b0011001111001100001100111100110001100110100110011001100101100110,
64'b1111111100000000111111110000000010101010101010101010101010101010,
64'b0101010110101010010101011010101001011010101001011010010101011010,
64'b1100110011001100110011001100110010100101101001010101101001011010,
64'b1100110000110011001100111100110010011001011001101001100101100110,
64'b0011001111001100001100111100110001010101010101011010101010101010,
64'b0101010110101010010101011010101010011001100110010110011001100110,
64'b1001011010010110100101101001011010100101010110101010010101011010,
64'b1001011010010110100101101001011000111100001111000011110000111100,
64'b1111000000001111000011111111000000110011001100111100110011001100,
64'b1111111100000000111111110000000000001111000011111111000011110000,
64'b1001011001101001011010011001011011111111111111110000000000000000,
64'b1100110011001100110011001100110001100110011001100110011001100110,
64'b0101101001011010010110100101101001101001011010011001011010010110,
64'b1001100101100110100110010110011001100110011001100110011001100110,
64'b0011001100110011110011001100110001100110100110011001100101100110,
64'b1111000011110000111100001111000010011001011001101001100101100110,
64'b0000111100001111111100001111000001101001011010011001011010010110,
64'b1010010110100101010110100101101011001100110011001100110011001100,
64'b0011001100110011110011001100110010010110100101101001011010010110,
64'b1100001100111100110000110011110001100110100110011001100101100110,
64'b1100001100111100110000110011110000001111111100000000111111110000,
64'b0000000011111111111111110000000011110000111100001111000011110000,
64'b0101010101010101101010101010101001010101101010100101010110101010,
64'b0011110011000011110000110011110010101010101010101010101010101010,
64'b0101101001011010010110100101101010010110100101101001011010010110,
64'b0011001111001100001100111100110011000011001111001100001100111100,
64'b0011110000111100001111000011110010010110100101101001011010010110,
64'b1111000011110000111100001111000011000011110000110011110000111100,
64'b0101010110101010010101011010101001101001011010011001011010010110,
64'b1111111100000000111111110000000011000011001111001100001100111100,
64'b1001100101100110100110010110011001011010010110100101101001011010,
64'b0101101001011010010110100101101011000011001111001100001100111100,
64'b0101101010100101101001010101101011000011110000110011110000111100,
64'b1111000000001111000011111111000010101010010101010101010110101010,
64'b1111111111111111000000000000000011111111000000001111111100000000,
64'b0110011001100110011001100110011000110011001100111100110011001100,
64'b0101101010100101101001010101101011001100110011001100110011001100,
64'b1001100101100110100110010110011011000011001111001100001100111100,
64'b0000111100001111111100001111000011110000000011110000111111110000,
64'b0000111111110000000011111111000011000011001111001100001100111100,
64'b0101010110101010010101011010101010100101010110101010010101011010,
64'b0011001100110011110011001100110001101001100101100110100110010110,
64'b1111111111111111000000000000000001011010101001011010010101011010,
64'b1100001111000011001111000011110000110011110011000011001111001100,
64'b0011001111001100001100111100110011110000000011110000111111110000,
64'b1100110000110011001100111100110000001111111100000000111111110000,
64'b1010101001010101010101011010101010011001100110010110011001100110,
64'b1010101010101010101010101010101001010101010101011010101010101010,
64'b1001011010010110100101101001011011110000111100001111000011110000,
64'b1100110000110011001100111100110001011010010110100101101001011010,
64'b0110100101101001100101101001011011110000000011110000111111110000,
64'b1111111100000000111111110000000000000000111111111111111100000000,
64'b0101010110101010010101011010101010100101010110101010010101011010,
64'b0110011001100110011001100110011011111111000000001111111100000000,
64'b0101010110101010010101011010101001011010101001011010010101011010,
64'b1111000011110000111100001111000001010101101010100101010110101010,
64'b0000111100001111111100001111000010010110011010010110100110010110,
64'b0000111100001111111100001111000010010110100101101001011010010110,
64'b1111000011110000111100001111000000110011110011000011001111001100,
64'b0101010110101010010101011010101000001111000011111111000011110000,
64'b1001100101100110100110010110011010011001100110010110011001100110,
64'b1001011001101001011010011001011011111111111111110000000000000000,
64'b1111111100000000111111110000000001011010101001011010010101011010,
64'b0011110000111100001111000011110000000000111111111111111100000000,
64'b1010101010101010101010101010101000110011001100111100110011001100,
64'b0000111111110000000011111111000010100101010110101010010101011010,
64'b1111000011110000111100001111000001010101010101011010101010101010,
64'b0110011010011001100110010110011011001100001100110011001111001100,
64'b0000111111110000000011111111000010011001100110010110011001100110,
64'b1111000000001111000011111111000000111100110000111100001100111100,
64'b0101101010100101101001010101101001101001100101100110100110010110,
64'b1010010101011010101001010101101000001111000011111111000011110000,
64'b0110011010011001100110010110011011111111000000001111111100000000,
64'b0101101010100101101001010101101010010110100101101001011010010110,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b1010101001010101010101011010101001100110100110011001100101100110,
64'b0011001111001100001100111100110001010101010101011010101010101010,
64'b0110011001100110011001100110011001011010010110100101101001011010,
64'b1111000011110000111100001111000010011001011001101001100101100110,
64'b0011001111001100001100111100110011001100110011001100110011001100,
64'b1001011001101001011010011001011010100101101001010101101001011010,
64'b0101101010100101101001010101101010010110100101101001011010010110,
64'b0000111111110000000011111111000001011010101001011010010101011010,
64'b0110100110010110011010011001011010010110011010010110100110010110,
64'b1001011001101001011010011001011011111111000000001111111100000000,
64'b1001011001101001011010011001011001010101010101011010101010101010,
64'b1111111111111111000000000000000011000011001111001100001100111100,
64'b1111000000001111000011111111000011001100110011001100110011001100,
64'b1100110000110011001100111100110011000011110000110011110000111100,
64'b1001100110011001011001100110011001100110011001100110011001100110,
64'b1001011010010110100101101001011010011001011001101001100101100110,
64'b1111000011110000111100001111000000111100001111000011110000111100,
64'b0000111100001111111100001111000011110000111100001111000011110000,
64'b0011110011000011110000110011110000110011110011000011001111001100,
64'b0110011010011001100110010110011001101001100101100110100110010110,
64'b1010101001010101010101011010101011001100001100110011001111001100,
64'b0011110011000011110000110011110010010110011010010110100110010110,
64'b0011110011000011110000110011110001010101010101011010101010101010,
64'b1001011001101001011010011001011011001100110011001100110011001100,
64'b1010101010101010101010101010101001011010101001011010010101011010,
64'b1010101001010101010101011010101011110000111100001111000011110000,
64'b1010010110100101010110100101101000001111111100000000111111110000,
64'b1001011010010110100101101001011010010110100101101001011010010110,
64'b0110100110010110011010011001011011000011110000110011110000111100,
64'b1111111100000000111111110000000000001111111100000000111111110000,
64'b1001100101100110100110010110011001010101101010100101010110101010,
64'b0000111100001111111100001111000000001111000011111111000011110000,
64'b1001100110011001011001100110011000111100110000111100001100111100,
64'b1001011010010110100101101001011000001111000011111111000011110000,
64'b0101010110101010010101011010101010010110011010010110100110010110,
64'b1010101001010101010101011010101001100110011001100110011001100110,
64'b1100001111000011001111000011110001011010010110100101101001011010,
64'b1111111100000000111111110000000011001100001100110011001111001100,
64'b1010010101011010101001010101101001010101101010100101010110101010,
64'b0110011001100110011001100110011000000000111111111111111100000000,
64'b0101010110101010010101011010101011000011001111001100001100111100,
64'b1001011001101001011010011001011000001111111100000000111111110000,
64'b0000111111110000000011111111000001010101101010100101010110101010,
64'b1010010110100101010110100101101000110011001100111100110011001100,
64'b1010101010101010101010101010101011111111000000001111111100000000,
64'b0110011001100110011001100110011001011010101001011010010101011010,
64'b0110011010011001100110010110011001010101101010100101010110101010,
64'b0011110000111100001111000011110010010110011010010110100110010110,
64'b1100001111000011001111000011110010010110100101101001011010010110,
64'b1111000011110000111100001111000000110011110011000011001111001100,
64'b1100110000110011001100111100110000001111000011111111000011110000,
64'b0101101001011010010110100101101010011001100110010110011001100110,
64'b1100001100111100110000110011110011111111111111110000000000000000,
64'b0000111100001111111100001111000001011010101001011010010101011010,
64'b1001011001101001011010011001011000000000111111111111111100000000,
64'b0101101001011010010110100101101011001100110011001100110011001100,
64'b1001100101100110100110010110011010010110100101101001011010010110,
64'b0110011001100110011001100110011000000000111111111111111100000000,
64'b0011110000111100001111000011110000111100110000111100001100111100,
64'b1100001111000011001111000011110010010110100101101001011010010110,
64'b1010010101011010101001010101101000110011110011000011001111001100,
64'b0000111111110000000011111111000010011001011001101001100101100110,
64'b0101010110101010010101011010101001011010101001011010010101011010,
64'b0000111100001111111100001111000001100110011001100110011001100110,
64'b1001100101100110100110010110011000000000111111111111111100000000,
64'b1111000000001111000011111111000001010101101010100101010110101010,
64'b1111111100000000111111110000000001011010101001011010010101011010,
64'b1001011001101001011010011001011011111111111111110000000000000000,
64'b1001100101100110100110010110011001010101101010100101010110101010,
64'b1010010110100101010110100101101000001111111100000000111111110000,
64'b0110100110010110011010011001011010101010010101010101010110101010,
64'b1111111100000000111111110000000010101010010101010101010110101010,
64'b0000000011111111111111110000000001100110100110011001100101100110,
64'b0110100110010110011010011001011000000000000000000000000000000000,
64'b1111000000001111000011111111000000110011001100111100110011001100,
64'b0110011010011001100110010110011010011001100110010110011001100110,
64'b0110011001100110011001100110011000001111111100000000111111110000,
64'b1111111100000000111111110000000001101001100101100110100110010110,
64'b1111111111111111000000000000000001100110100110011001100101100110,
64'b0110100101101001100101101001011011110000000011110000111111110000,
64'b1001011001101001011010011001011000000000000000000000000000000000,
64'b1001100101100110100110010110011001101001100101100110100110010110,
64'b1111111100000000111111110000000010101010010101010101010110101010,
64'b1100001111000011001111000011110000110011001100111100110011001100,
64'b0000111100001111111100001111000010011001100110010110011001100110,
64'b1111000011110000111100001111000001101001011010011001011010010110,
64'b1001100101100110100110010110011010101010101010101010101010101010,
64'b1111000000001111000011111111000011110000111100001111000011110000,
64'b0011110011000011110000110011110010010110100101101001011010010110,
64'b0000111111110000000011111111000010101010010101010101010110101010,
64'b0110100110010110011010011001011000111100110000111100001100111100,
64'b1111111100000000111111110000000011000011110000110011110000111100,
64'b0101010110101010010101011010101010101010010101010101010110101010,
64'b0011110011000011110000110011110010101010101010101010101010101010,
64'b1001100101100110100110010110011011000011001111001100001100111100,
64'b1111111111111111000000000000000010011001100110010110011001100110,
64'b0000111111110000000011111111000001011010010110100101101001011010,
64'b0101010110101010010101011010101010010110100101101001011010010110,
64'b0101010110101010010101011010101001101001100101100110100110010110,
64'b1100001111000011001111000011110001100110011001100110011001100110,
64'b0000000011111111111111110000000011111111000000001111111100000000,
64'b0101101010100101101001010101101011000011001111001100001100111100,
64'b1010101001010101010101011010101000110011001100111100110011001100,
64'b0011110011000011110000110011110001011010101001011010010101011010,
64'b1111111111111111000000000000000010100101010110101010010101011010,
64'b0011001100110011110011001100110010011001100110010110011001100110,
64'b1111000000001111000011111111000001100110011001100110011001100110,
64'b1001011010010110100101101001011000001111111100000000111111110000,
64'b0110011001100110011001100110011011110000111100001111000011110000,
64'b1111111111111111000000000000000011001100110011001100110011001100,
64'b1100001111000011001111000011110000110011110011000011001111001100,
64'b0011110000111100001111000011110000110011110011000011001111001100,
64'b0000000011111111111111110000000000110011001100111100110011001100,
64'b1010010110100101010110100101101000001111000011111111000011110000,
64'b0011001100110011110011001100110010100101101001010101101001011010,
64'b0000000011111111111111110000000001101001100101100110100110010110,
64'b1100110011001100110011001100110011110000111100001111000011110000,
64'b0101010110101010010101011010101010011001100110010110011001100110,
64'b0110011001100110011001100110011000000000000000000000000000000000,
64'b0000000011111111111111110000000000111100001111000011110000111100,
64'b0110011001100110011001100110011011110000111100001111000011110000,
64'b0101101001011010010110100101101001010101101010100101010110101010,
64'b0101010110101010010101011010101011110000111100001111000011110000,
64'b0101010110101010010101011010101000001111000011111111000011110000,
64'b1010101001010101010101011010101000001111000011111111000011110000,
64'b1111000011110000111100001111000011110000111100001111000011110000,
64'b0110100110010110011010011001011001010101101010100101010110101010,
64'b0000111111110000000011111111000010011001011001101001100101100110,
64'b1100110000110011001100111100110010010110011010010110100110010110,
64'b1100110000110011001100111100110011111111000000001111111100000000,
64'b1100110000110011001100111100110000111100001111000011110000111100,
64'b0000000000000000000000000000000010101010101010101010101010101010,
64'b0101010101010101101010101010101000001111111100000000111111110000,
64'b1001100101100110100110010110011011111111000000001111111100000000,
64'b1111111100000000111111110000000000110011001100111100110011001100,
64'b0110011010011001100110010110011011111111000000001111111100000000,
64'b1100001111000011001111000011110011111111000000001111111100000000,
64'b0011110000111100001111000011110001010101101010100101010110101010,
64'b0101101010100101101001010101101001010101101010100101010110101010,
64'b1100110000110011001100111100110000110011001100111100110011001100,
64'b0101010101010101101010101010101011000011110000110011110000111100,
64'b1001011001101001011010011001011000111100110000111100001100111100,
64'b0011001111001100001100111100110001010101010101011010101010101010,
64'b0101101010100101101001010101101000001111111100000000111111110000,
64'b1001011010010110100101101001011011001100110011001100110011001100,
64'b0110011001100110011001100110011000000000111111111111111100000000,
64'b1001100101100110100110010110011000000000000000000000000000000000,
64'b0101010101010101101010101010101011110000111100001111000011110000,
64'b1100001111000011001111000011110001010101010101011010101010101010,
64'b1010010101011010101001010101101011111111111111110000000000000000,
64'b1010010101011010101001010101101000110011001100111100110011001100,
64'b1100110000110011001100111100110000110011001100111100110011001100,
64'b1010010110100101010110100101101011110000111100001111000011110000,
64'b0110011001100110011001100110011010100101010110101010010101011010,
64'b1001011001101001011010011001011001011010101001011010010101011010,
64'b1010010110100101010110100101101001100110011001100110011001100110,
64'b1100110000110011001100111100110010101010010101010101010110101010,
64'b0110100110010110011010011001011011110000111100001111000011110000,
64'b0011110000111100001111000011110011111111111111110000000000000000,
64'b0011110000111100001111000011110010101010101010101010101010101010,
64'b1100110011001100110011001100110011111111000000001111111100000000,
64'b1010010101011010101001010101101011001100110011001100110011001100,
64'b0110011010011001100110010110011010101010101010101010101010101010,
64'b1100110000110011001100111100110001011010010110100101101001011010,
64'b0000111100001111111100001111000001011010010110100101101001011010,
64'b1001100101100110100110010110011001010101101010100101010110101010,
64'b1001011010010110100101101001011011001100001100110011001111001100,
64'b0011110011000011110000110011110011001100001100110011001111001100,
64'b1001100101100110100110010110011010010110100101101001011010010110,
64'b1010010110100101010110100101101000110011001100111100110011001100,
64'b1001011001101001011010011001011001010101101010100101010110101010,
64'b0000111111110000000011111111000000000000000000000000000000000000,
64'b0000111111110000000011111111000001100110011001100110011001100110,
64'b0101101001011010010110100101101001010101010101011010101010101010,
64'b1100110000110011001100111100110011110000111100001111000011110000,
64'b1100001111000011001111000011110011001100110011001100110011001100,
64'b1010010110100101010110100101101000110011110011000011001111001100,
64'b0101010110101010010101011010101000110011110011000011001111001100,
64'b0110100101101001100101101001011000110011001100111100110011001100,
64'b1100001100111100110000110011110000001111000011111111000011110000,
64'b1111000000001111000011111111000010100101101001010101101001011010,
64'b0110100101101001100101101001011001101001100101100110100110010110,
64'b0011001111001100001100111100110011110000111100001111000011110000,
64'b1001011001101001011010011001011010011001100110010110011001100110,
64'b1010101001010101010101011010101000000000000000000000000000000000,
64'b1111111100000000111111110000000000111100001111000011110000111100,
64'b1111111111111111000000000000000010011001011001101001100101100110,
64'b0011110011000011110000110011110011001100001100110011001111001100,
64'b1001100110011001011001100110011010100101101001010101101001011010,
64'b0101010101010101101010101010101011001100110011001100110011001100,
64'b0101101010100101101001010101101011000011110000110011110000111100,
64'b1010101001010101010101011010101001011010101001011010010101011010,
64'b1010010110100101010110100101101010100101101001010101101001011010,
64'b1100110011001100110011001100110011111111000000001111111100000000,
64'b1010101010101010101010101010101011001100110011001100110011001100,
64'b1100110000110011001100111100110001100110100110011001100101100110,
64'b1111000011110000111100001111000010010110100101101001011010010110,
64'b1100110000110011001100111100110010101010101010101010101010101010,
64'b1111000011110000111100001111000010100101010110101010010101011010,
64'b0101010101010101101010101010101001101001011010011001011010010110,
64'b0110011001100110011001100110011000001111000011111111000011110000,
64'b0000111100001111111100001111000010011001011001101001100101100110,
64'b0011001100110011110011001100110001011010010110100101101001011010,
64'b0011110000111100001111000011110000001111111100000000111111110000,
64'b0011001111001100001100111100110001100110100110011001100101100110,
64'b0011110011000011110000110011110010011001011001101001100101100110,
64'b1001011010010110100101101001011001010101010101011010101010101010,
64'b0110011001100110011001100110011011110000111100001111000011110000,
64'b1100001100111100110000110011110011000011110000110011110000111100,
64'b1010010101011010101001010101101001101001100101100110100110010110,
64'b1100001100111100110000110011110011001100110011001100110011001100,
64'b1010010101011010101001010101101000110011110011000011001111001100,
64'b0011001100110011110011001100110001101001100101100110100110010110,
64'b1010101001010101010101011010101001010101101010100101010110101010,
64'b0110011010011001100110010110011001101001011010011001011010010110,
64'b0000111100001111111100001111000000110011110011000011001111001100,
64'b1111111111111111000000000000000000000000111111111111111100000000,
64'b1010010101011010101001010101101011000011110000110011110000111100,
64'b0101010110101010010101011010101001101001011010011001011010010110,
64'b1010010101011010101001010101101011001100110011001100110011001100,
64'b1001011010010110100101101001011001010101101010100101010110101010,
64'b0011110000111100001111000011110000001111111100000000111111110000,
64'b0011110011000011110000110011110010010110011010010110100110010110,
64'b0011110000111100001111000011110011110000111100001111000011110000,
64'b1100001100111100110000110011110011110000111100001111000011110000,
64'b1111000011110000111100001111000000111100110000111100001100111100,
64'b1001100110011001011001100110011000110011001100111100110011001100,
64'b0110100101101001100101101001011011000011001111001100001100111100,
64'b0101010110101010010101011010101010100101101001010101101001011010,
64'b1010101010101010101010101010101011111111111111110000000000000000,
64'b0110011010011001100110010110011010100101010110101010010101011010,
64'b0011001100110011110011001100110001101001100101100110100110010110,
64'b1100110000110011001100111100110001011010010110100101101001011010,
64'b1100001100111100110000110011110000110011001100111100110011001100,
64'b0000111111110000000011111111000000000000111111111111111100000000,
64'b1111000000001111000011111111000000111100110000111100001100111100,
64'b1010010101011010101001010101101001010101101010100101010110101010,
64'b0000111111110000000011111111000011111111000000001111111100000000,
64'b1010101001010101010101011010101001011010101001011010010101011010,
64'b0000000011111111111111110000000001011010010110100101101001011010,
64'b1111000000001111000011111111000001011010101001011010010101011010,
64'b1100110011001100110011001100110000110011110011000011001111001100,
64'b1001011001101001011010011001011010101010101010101010101010101010,
64'b0110100110010110011010011001011001100110100110011001100101100110,
64'b1111111111111111000000000000000000111100110000111100001100111100,
64'b0110100101101001100101101001011000110011110011000011001111001100,
64'b1111000000001111000011111111000011110000111100001111000011110000,
64'b1100110011001100110011001100110001010101010101011010101010101010,
64'b1111000000001111000011111111000001011010101001011010010101011010,
64'b1010101010101010101010101010101010011001100110010110011001100110,
64'b0000111111110000000011111111000000000000000000000000000000000000,
64'b0110011001100110011001100110011001100110100110011001100101100110,
64'b0110100110010110011010011001011010011001011001101001100101100110,
64'b0011001111001100001100111100110011001100001100110011001111001100,
64'b0000111100001111111100001111000010100101101001010101101001011010,
64'b0110011001100110011001100110011011001100110011001100110011001100,
64'b0011110000111100001111000011110011000011110000110011110000111100,
64'b1010010110100101010110100101101001011010101001011010010101011010,
64'b1010010101011010101001010101101010100101101001010101101001011010,
64'b0000000011111111111111110000000011111111000000001111111100000000,
64'b1001011001101001011010011001011011001100110011001100110011001100,
64'b1111000000001111000011111111000001100110100110011001100101100110,
64'b1010101001010101010101011010101010010110100101101001011010010110,
64'b0000111111110000000011111111000010101010101010101010101010101010,
64'b0011110000111100001111000011110000111100001111000011110000111100,
64'b0011110011000011110000110011110001010101101010100101010110101010,
64'b0000111100001111111100001111000010010110100101101001011010010110,
64'b1111111100000000111111110000000011001100001100110011001111001100,
64'b1001011010010110100101101001011000000000111111111111111100000000,
64'b0000111111110000000011111111000010100101101001010101101001011010,
64'b0011001111001100001100111100110011000011001111001100001100111100,
64'b0110011010011001100110010110011001010101101010100101010110101010,
64'b1111111111111111000000000000000011111111111111110000000000000000,
64'b1001011001101001011010011001011000111100110000111100001100111100,
64'b1010101001010101010101011010101000110011001100111100110011001100,
64'b1001100110011001011001100110011010100101101001010101101001011010,
64'b0101010110101010010101011010101000111100001111000011110000111100,
64'b0101101010100101101001010101101001011010101001011010010101011010,
64'b1100110011001100110011001100110000001111111100000000111111110000,
64'b1100110000110011001100111100110001011010101001011010010101011010,
64'b0000000000000000000000000000000001011010010110100101101001011010,
64'b1001100110011001011001100110011000001111111100000000111111110000,
64'b1010101010101010101010101010101000110011001100111100110011001100,
64'b1010101010101010101010101010101011111111000000001111111100000000,
64'b0000111100001111111100001111000011111111111111110000000000000000,
64'b0000000000000000000000000000000010101010101010101010101010101010,
64'b0101101001011010010110100101101010010110100101101001011010010110,
64'b0110100101101001100101101001011010101010101010101010101010101010,
64'b0101101010100101101001010101101001010101010101011010101010101010,
64'b1001011010010110100101101001011001010101101010100101010110101010,
64'b1001100101100110100110010110011001100110100110011001100101100110,
64'b0110011010011001100110010110011010101010010101010101010110101010,
64'b1001011010010110100101101001011011001100001100110011001111001100,
64'b1111111111111111000000000000000010011001011001101001100101100110,
64'b0110011010011001100110010110011000000000111111111111111100000000,
64'b1100110000110011001100111100110011110000111100001111000011110000,
64'b0110100101101001100101101001011001010101010101011010101010101010,
64'b0011001111001100001100111100110000000000000000000000000000000000,
64'b0000000000000000000000000000000001100110011001100110011001100110,
64'b1111111111111111000000000000000011000011001111001100001100111100,
64'b0011001111001100001100111100110011001100110011001100110011001100,
64'b1010101010101010101010101010101011001100110011001100110011001100,
64'b1001100101100110100110010110011001100110011001100110011001100110,
64'b0110100101101001100101101001011001101001011010011001011010010110,
64'b1100001111000011001111000011110010011001100110010110011001100110,
64'b0110100110010110011010011001011010100101101001010101101001011010,
64'b0000000000000000000000000000000001101001011010011001011010010110,
64'b0110100101101001100101101001011011111111111111110000000000000000,
64'b1010010110100101010110100101101001010101101010100101010110101010,
64'b0110100110010110011010011001011011001100110011001100110011001100,
64'b1010010110100101010110100101101010101010101010101010101010101010,
64'b0000000000000000000000000000000000111100001111000011110000111100,
64'b0000000000000000000000000000000011110000000011110000111111110000,
64'b1010010110100101010110100101101011110000111100001111000011110000,
64'b1100110011001100110011001100110011110000111100001111000011110000,
64'b0011110000111100001111000011110000111100001111000011110000111100,
64'b0011110011000011110000110011110010010110011010010110100110010110,
64'b1001100110011001011001100110011010101010010101010101010110101010,
64'b0000111111110000000011111111000000000000111111111111111100000000,
64'b0101010101010101101010101010101000111100110000111100001100111100,
64'b1001100110011001011001100110011011110000000011110000111111110000,
64'b0011001100110011110011001100110000110011110011000011001111001100,
64'b0011001111001100001100111100110001010101010101011010101010101010,
64'b1111111100000000111111110000000000000000000000000000000000000000,
64'b0000000000000000000000000000000010100101010110101010010101011010,
64'b1100110000110011001100111100110011001100110011001100110011001100,
64'b1100001100111100110000110011110010100101010110101010010101011010,
64'b1001011001101001011010011001011000110011001100111100110011001100,
64'b1111111100000000111111110000000011111111000000001111111100000000,
64'b0000111111110000000011111111000000111100110000111100001100111100,
64'b1010101001010101010101011010101010011001100110010110011001100110,
64'b0011001111001100001100111100110001010101010101011010101010101010,
64'b1001100110011001011001100110011001011010101001011010010101011010,
64'b1100110000110011001100111100110010101010010101010101010110101010,
64'b1111000000001111000011111111000010100101101001010101101001011010,
64'b0000000000000000000000000000000011001100110011001100110011001100,
64'b0011001100110011110011001100110010101010101010101010101010101010,
64'b1010101010101010101010101010101011001100001100110011001111001100,
64'b1100001100111100110000110011110011110000111100001111000011110000,
64'b1010101001010101010101011010101011001100001100110011001111001100,
64'b1111000011110000111100001111000011110000111100001111000011110000,
64'b0101101001011010010110100101101010101010101010101010101010101010,
64'b0101010110101010010101011010101001011010101001011010010101011010,
64'b0000111111110000000011111111000010010110100101101001011010010110,
64'b0011110000111100001111000011110001100110011001100110011001100110,
64'b0110100101101001100101101001011001100110100110011001100101100110,
64'b1111111100000000111111110000000010011001100110010110011001100110,
64'b0000000000000000000000000000000010011001011001101001100101100110,
64'b0000111100001111111100001111000001011010010110100101101001011010,
64'b0011110000111100001111000011110011001100110011001100110011001100,
64'b1100110011001100110011001100110000001111000011111111000011110000,
64'b0011110000111100001111000011110001010101101010100101010110101010,
64'b1100001111000011001111000011110000001111000011111111000011110000,
64'b1001100110011001011001100110011001010101101010100101010110101010,
64'b1100001100111100110000110011110011001100110011001100110011001100,
64'b1001100110011001011001100110011011001100001100110011001111001100,
64'b0000000011111111111111110000000001101001100101100110100110010110,
64'b0000111111110000000011111111000000111100001111000011110000111100,
64'b1100001100111100110000110011110011000011110000110011110000111100,
64'b0101010101010101101010101010101010010110100101101001011010010110,
64'b0000000000000000000000000000000001101001011010011001011010010110,
64'b1111111100000000111111110000000000110011110011000011001111001100,
64'b1010010101011010101001010101101011110000111100001111000011110000,
64'b1111000011110000111100001111000011111111000000001111111100000000,
64'b0000111111110000000011111111000010011001100110010110011001100110,
64'b0000111111110000000011111111000011111111000000001111111100000000,
64'b1001011010010110100101101001011010011001100110010110011001100110,
64'b1010010101011010101001010101101011110000111100001111000011110000,
64'b0011110000111100001111000011110000001111000011111111000011110000,
64'b0101010101010101101010101010101010010110011010010110100110010110,
64'b1010101001010101010101011010101000001111111100000000111111110000,
64'b1111000000001111000011111111000000001111111100000000111111110000,
64'b1100110011001100110011001100110001101001100101100110100110010110,
64'b1010101010101010101010101010101011000011001111001100001100111100,
64'b1111111111111111000000000000000010100101101001010101101001011010,
64'b1100110000110011001100111100110011111111000000001111111100000000,
64'b1111111100000000111111110000000011111111111111110000000000000000,
64'b0000000011111111111111110000000000111100001111000011110000111100,
64'b0000000011111111111111110000000001010101010101011010101010101010,
64'b1100001100111100110000110011110000111100001111000011110000111100,
64'b0011001111001100001100111100110001010101101010100101010110101010,
64'b1010010101011010101001010101101011111111000000001111111100000000,
64'b1100110011001100110011001100110010010110011010010110100110010110,
64'b1001100110011001011001100110011010101010010101010101010110101010,
64'b1010101001010101010101011010101000000000111111111111111100000000,
64'b0101101001011010010110100101101000111100110000111100001100111100,
64'b1100110011001100110011001100110011110000000011110000111111110000,
64'b0000000000000000000000000000000000110011110011000011001111001100,
64'b1010010110100101010110100101101001010101010101011010101010101010,
64'b0101010101010101101010101010101000000000000000000000000000000000,
64'b1111111111111111000000000000000010100101010110101010010101011010,
64'b0101010101010101101010101010101011001100110011001100110011001100,
64'b0101101010100101101001010101101010100101010110101010010101011010,
64'b1111000011110000111100001111000011001100110011001100110011001100,
64'b1100110011001100110011001100110000001111111100000000111111110000,
64'b1010010101011010101001010101101010010110011010010110100110010110,
64'b0101101010100101101001010101101011000011110000110011110000111100,
64'b0000000011111111111111110000000010100101101001010101101001011010,
64'b1111000000001111000011111111000000111100110000111100001100111100,
64'b0000000000000000000000000000000011001100001100110011001111001100,
64'b0000000011111111111111110000000010010110011010010110100110010110,
64'b1010010101011010101001010101101011111111111111110000000000000000,
64'b0011001111001100001100111100110010101010010101010101010110101010,
64'b0000000000000000000000000000000011000011110000110011110000111100,
64'b1100001100111100110000110011110011110000111100001111000011110000,
64'b0110100110010110011010011001011000000000000000000000000000000000,
64'b0011001111001100001100111100110011110000111100001111000011110000,
64'b0011110000111100001111000011110010101010010101010101010110101010,
64'b0110100101101001100101101001011000111100110000111100001100111100,
64'b1001011010010110100101101001011010100101010110101010010101011010,
64'b0101010110101010010101011010101010011001011001101001100101100110,
64'b0101101001011010010110100101101001011010101001011010010101011010,
64'b1010101010101010101010101010101010100101101001010101101001011010,
64'b1111111100000000111111110000000010010110011010010110100110010110,
64'b1100001111000011001111000011110010101010101010101010101010101010,
64'b0011110011000011110000110011110010011001100110010110011001100110,
64'b0000000000000000000000000000000010100101010110101010010101011010,
64'b0011001100110011110011001100110001010101101010100101010110101010,
64'b0101010101010101101010101010101000000000000000000000000000000000,
64'b1100001100111100110000110011110011111111000000001111111100000000,
64'b0110100110010110011010011001011010011001100110010110011001100110,
64'b0110011001100110011001100110011001011010101001011010010101011010,
64'b0011001100110011110011001100110001100110100110011001100101100110,
64'b0011001111001100001100111100110011000011110000110011110000111100,
64'b1100001111000011001111000011110011001100001100110011001111001100,
64'b1100110011001100110011001100110010011001011001101001100101100110,
64'b1111111100000000111111110000000010010110011010010110100110010110,
64'b1010101010101010101010101010101001100110011001100110011001100110,
64'b0110100101101001100101101001011000111100001111000011110000111100,
64'b1010101010101010101010101010101001100110100110011001100101100110,
64'b0011001111001100001100111100110000110011001100111100110011001100,
64'b0000111111110000000011111111000000000000000000000000000000000000,
64'b1001011010010110100101101001011000000000000000000000000000000000,
64'b1001011001101001011010011001011000111100001111000011110000111100,
64'b0011110000111100001111000011110001100110100110011001100101100110,
64'b1111000011110000111100001111000001101001011010011001011010010110,
64'b1010010110100101010110100101101010100101010110101010010101011010,
64'b0000111111110000000011111111000010100101101001010101101001011010,
64'b0101101001011010010110100101101001101001011010011001011010010110,
64'b1111111111111111000000000000000000111100110000111100001100111100,
64'b1100110011001100110011001100110010010110100101101001011010010110,
64'b1100001100111100110000110011110000001111111100000000111111110000,
64'b0110011001100110011001100110011011000011110000110011110000111100,
64'b0000111100001111111100001111000001011010010110100101101001011010,
64'b0000000011111111111111110000000010101010101010101010101010101010,
64'b1100001100111100110000110011110000000000000000000000000000000000,
64'b0101101010100101101001010101101010100101010110101010010101011010,
64'b0000000000000000000000000000000011000011110000110011110000111100,
64'b1010010110100101010110100101101001101001100101100110100110010110,
64'b0011001100110011110011001100110001100110100110011001100101100110,
64'b0101101001011010010110100101101000110011110011000011001111001100,
64'b0011001111001100001100111100110001101001100101100110100110010110,
64'b0000000011111111111111110000000001011010101001011010010101011010,
64'b1111111100000000111111110000000001101001100101100110100110010110,
64'b1100001111000011001111000011110000000000111111111111111100000000,
64'b0011110000111100001111000011110000001111111100000000111111110000,
64'b0011110000111100001111000011110010011001011001101001100101100110,
64'b0011110011000011110000110011110011001100110011001100110011001100,
64'b1001011010010110100101101001011000000000000000000000000000000000,
64'b1010101001010101010101011010101011001100001100110011001111001100,
64'b0000111111110000000011111111000000001111111100000000111111110000,
64'b0110100101101001100101101001011010010110011010010110100110010110,
64'b0101101010100101101001010101101011000011110000110011110000111100,
64'b0110100101101001100101101001011010100101101001010101101001011010,
64'b0000111100001111111100001111000000111100110000111100001100111100,
64'b1111111100000000111111110000000011001100001100110011001111001100,
64'b1111000000001111000011111111000010010110011010010110100110010110,
64'b0011110000111100001111000011110011111111111111110000000000000000,
64'b1010010101011010101001010101101010101010010101010101010110101010,
64'b1100110011001100110011001100110011000011110000110011110000111100,
64'b1001100110011001011001100110011011110000111100001111000011110000,
64'b0101101001011010010110100101101000000000000000000000000000000000,
64'b1001100110011001011001100110011011000011110000110011110000111100,
64'b1010101001010101010101011010101000001111000011111111000011110000,
64'b1100001100111100110000110011110001100110011001100110011001100110,
64'b0110011010011001100110010110011010100101101001010101101001011010,
64'b0110100110010110011010011001011001101001011010011001011010010110,
64'b0101010110101010010101011010101001011010101001011010010101011010,
64'b0101010101010101101010101010101010100101010110101010010101011010,
64'b0000000011111111111111110000000000110011001100111100110011001100,
64'b1010010101011010101001010101101010011001011001101001100101100110,
64'b1100110000110011001100111100110010011001100110010110011001100110,
64'b1111000011110000111100001111000001100110011001100110011001100110,
64'b0011110000111100001111000011110000111100001111000011110000111100,
64'b1001100101100110100110010110011000110011110011000011001111001100,
64'b0101101001011010010110100101101011000011001111001100001100111100,
64'b0011110011000011110000110011110011110000111100001111000011110000,
64'b0000000000000000000000000000000011001100001100110011001111001100,
64'b1100001100111100110000110011110000110011001100111100110011001100,
64'b0110011001100110011001100110011010011001100110010110011001100110,
64'b0011001100110011110011001100110001100110100110011001100101100110,
64'b1100110000110011001100111100110001100110011001100110011001100110,
64'b1111000000001111000011111111000001010101101010100101010110101010,
64'b0101010101010101101010101010101001011010101001011010010101011010,
64'b0000111100001111111100001111000000111100001111000011110000111100,
64'b1001011010010110100101101001011001010101101010100101010110101010,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b0000111111110000000011111111000011000011001111001100001100111100,
64'b1111111100000000111111110000000001011010101001011010010101011010,
64'b0101010101010101101010101010101011111111000000001111111100000000,
64'b1111000000001111000011111111000000001111000011111111000011110000,
64'b1111000011110000111100001111000001011010010110100101101001011010,
64'b1100110000110011001100111100110010010110100101101001011010010110,
64'b1111000011110000111100001111000001101001011010011001011010010110,
64'b1010010101011010101001010101101010010110100101101001011010010110,
64'b0000111100001111111100001111000000110011001100111100110011001100,
64'b0101010110101010010101011010101011001100001100110011001111001100,
64'b0101010110101010010101011010101010100101010110101010010101011010,
64'b1010101010101010101010101010101000110011001100111100110011001100,
64'b0101010110101010010101011010101000111100001111000011110000111100,
64'b1100110011001100110011001100110000001111111100000000111111110000,
64'b0101010101010101101010101010101011001100001100110011001111001100,
64'b1100110011001100110011001100110001010101010101011010101010101010,
64'b1010101001010101010101011010101011111111000000001111111100000000,
64'b0101010110101010010101011010101010011001011001101001100101100110,
64'b0000111100001111111100001111000011000011001111001100001100111100,
64'b0101010110101010010101011010101011000011001111001100001100111100,
64'b1100110000110011001100111100110001101001100101100110100110010110,
64'b1111111100000000111111110000000011110000111100001111000011110000,
64'b1001100110011001011001100110011010100101101001010101101001011010,
64'b0011001100110011110011001100110001100110100110011001100101100110,
64'b1100110011001100110011001100110011110000111100001111000011110000,
64'b0011001100110011110011001100110010100101010110101010010101011010,
64'b1111000011110000111100001111000011111111000000001111111100000000,
64'b0000000000000000000000000000000011000011110000110011110000111100,
64'b1111111100000000111111110000000011000011001111001100001100111100,
64'b0110100110010110011010011001011000001111111100000000111111110000,
64'b1001100101100110100110010110011011000011001111001100001100111100,
64'b0000111100001111111100001111000000000000000000000000000000000000,
64'b1001100110011001011001100110011011110000000011110000111111110000,
64'b0000111111110000000011111111000000111100001111000011110000111100,
64'b1111000000001111000011111111000001011010010110100101101001011010,
64'b0000111111110000000011111111000000000000000000000000000000000000,
64'b0101101001011010010110100101101001101001011010011001011010010110,
64'b1001100101100110100110010110011010010110100101101001011010010110,
64'b1001100101100110100110010110011010100101101001010101101001011010,
64'b0110011001100110011001100110011000110011110011000011001111001100,
64'b0110011001100110011001100110011010100101010110101010010101011010,
64'b0101101010100101101001010101101001011010101001011010010101011010,
64'b0110011001100110011001100110011000000000111111111111111100000000,
64'b1100001100111100110000110011110011110000000011110000111111110000,
64'b0000111100001111111100001111000000000000000000000000000000000000,
64'b1001011010010110100101101001011000000000111111111111111100000000,
64'b1010101010101010101010101010101010100101010110101010010101011010,
64'b1010010110100101010110100101101000110011110011000011001111001100,
64'b1001100110011001011001100110011000000000000000000000000000000000,
64'b0011001111001100001100111100110011000011001111001100001100111100,
64'b0000000011111111111111110000000001101001100101100110100110010110,
64'b1010101001010101010101011010101000110011110011000011001111001100,
64'b0000111111110000000011111111000001011010010110100101101001011010,
64'b1111000011110000111100001111000011001100001100110011001111001100,
64'b0110100101101001100101101001011011001100001100110011001111001100,
64'b1100110000110011001100111100110001010101010101011010101010101010,
64'b1111000011110000111100001111000010101010010101010101010110101010,
64'b0000111100001111111100001111000010101010101010101010101010101010,
64'b0110100110010110011010011001011011111111111111110000000000000000,
64'b1100110000110011001100111100110001100110100110011001100101100110,
64'b1001011010010110100101101001011000001111000011111111000011110000,
64'b1010010101011010101001010101101000000000000000000000000000000000,
64'b1010010110100101010110100101101011110000000011110000111111110000,
64'b0011110011000011110000110011110000111100110000111100001100111100,
64'b1111000000001111000011111111000000001111000011111111000011110000,
64'b0110011001100110011001100110011000110011110011000011001111001100,
64'b0101010110101010010101011010101000001111000011111111000011110000,
64'b1100001100111100110000110011110010100101101001010101101001011010,
64'b1010010110100101010110100101101001100110011001100110011001100110,
64'b0101010110101010010101011010101010011001100110010110011001100110,
64'b1111111100000000111111110000000001100110011001100110011001100110,
64'b1001011001101001011010011001011000000000000000000000000000000000,
64'b0000111100001111111100001111000001101001011010011001011010010110,
64'b0110100110010110011010011001011001010101101010100101010110101010,
64'b1100110000110011001100111100110010101010101010101010101010101010,
64'b0011001111001100001100111100110000000000111111111111111100000000,
64'b0101101010100101101001010101101001011010101001011010010101011010,
64'b1010101001010101010101011010101001010101101010100101010110101010,
64'b1001011010010110100101101001011001011010010110100101101001011010,
64'b1001100110011001011001100110011011111111000000001111111100000000,
64'b1111000000001111000011111111000010011001011001101001100101100110,
64'b0011001111001100001100111100110010010110100101101001011010010110,
64'b1001100110011001011001100110011000111100001111000011110000111100,
64'b1111111111111111000000000000000010010110100101101001011010010110,
64'b0011110011000011110000110011110000000000000000000000000000000000,
64'b0101010110101010010101011010101011000011001111001100001100111100,
64'b1001011001101001011010011001011010011001100110010110011001100110,
64'b0000111100001111111100001111000011001100110011001100110011001100,
64'b1010010110100101010110100101101011111111111111110000000000000000,
64'b1100110000110011001100111100110001100110100110011001100101100110,
64'b1001100110011001011001100110011010011001100110010110011001100110,
64'b0110100110010110011010011001011000110011110011000011001111001100,
64'b1001011010010110100101101001011001010101010101011010101010101010,
64'b1010101001010101010101011010101011000011110000110011110000111100,
64'b1010010110100101010110100101101011000011001111001100001100111100,
64'b0011110000111100001111000011110000001111111100000000111111110000,
64'b1010101010101010101010101010101011000011001111001100001100111100,
64'b0101101010100101101001010101101000000000000000000000000000000000,
64'b1001100110011001011001100110011011110000000011110000111111110000,
64'b0011110011000011110000110011110000111100001111000011110000111100,
64'b0101010110101010010101011010101001011010010110100101101001011010,
64'b1001100101100110100110010110011000000000000000000000000000000000,
64'b1010010110100101010110100101101001101001011010011001011010010110,
64'b1001011010010110100101101001011010010110100101101001011010010110,
64'b0110100110010110011010011001011001011010010110100101101001011010,
64'b0011001111001100001100111100110010101010010101010101010110101010,
64'b1001100101100110100110010110011011111111000000001111111100000000,
64'b1010101001010101010101011010101011000011110000110011110000111100,
64'b0011110011000011110000110011110001101001011010011001011010010110,
64'b1010101001010101010101011010101000000000000000000000000000000000,
64'b0011110011000011110000110011110001010101101010100101010110101010,
64'b1001011010010110100101101001011001010101101010100101010110101010,
64'b0110100110010110011010011001011000001111000011111111000011110000,
64'b0000000011111111111111110000000011111111000000001111111100000000,
64'b0011001111001100001100111100110010011001100110010110011001100110,
64'b0101010110101010010101011010101000111100110000111100001100111100,
64'b1111000000001111000011111111000000111100001111000011110000111100,
64'b0110011001100110011001100110011011001100110011001100110011001100,
64'b1001011001101001011010011001011000110011001100111100110011001100,
64'b0101101010100101101001010101101001010101010101011010101010101010,
64'b1001100101100110100110010110011000001111111100000000111111110000,
64'b0110011001100110011001100110011001101001100101100110100110010110,
64'b0011001111001100001100111100110010101010101010101010101010101010,
64'b0110011001100110011001100110011000110011001100111100110011001100,
64'b1111111100000000111111110000000000110011001100111100110011001100,
64'b0101010101010101101010101010101011111111000000001111111100000000,
64'b1111111100000000111111110000000001010101010101011010101010101010,
64'b1001011001101001011010011001011000111100001111000011110000111100,
64'b0110011010011001100110010110011001011010101001011010010101011010,
64'b1111000011110000111100001111000010100101010110101010010101011010,
64'b1111000011110000111100001111000011110000111100001111000011110000,
64'b1010010110100101010110100101101001011010010110100101101001011010,
64'b1111111111111111000000000000000001100110011001100110011001100110,
64'b1100001100111100110000110011110010101010010101010101010110101010,
64'b0000000011111111111111110000000000111100110000111100001100111100,
64'b1010010101011010101001010101101011001100110011001100110011001100,
64'b0000000011111111111111110000000011110000111100001111000011110000,
64'b0110100101101001100101101001011001011010010110100101101001011010,
64'b1010010101011010101001010101101001010101010101011010101010101010,
64'b0101010110101010010101011010101011001100110011001100110011001100,
64'b0000111100001111111100001111000010100101010110101010010101011010,
64'b0011110011000011110000110011110011001100001100110011001111001100,
64'b1010010110100101010110100101101001100110100110011001100101100110,
64'b1001100101100110100110010110011011111111000000001111111100000000,
64'b0011001111001100001100111100110000110011110011000011001111001100,
64'b1010101010101010101010101010101000111100001111000011110000111100,
64'b0101101010100101101001010101101000110011001100111100110011001100,
64'b1111111111111111000000000000000001011010101001011010010101011010,
64'b0110011010011001100110010110011001011010010110100101101001011010,
64'b1111111111111111000000000000000011111111000000001111111100000000,
64'b0110100110010110011010011001011000110011110011000011001111001100,
64'b0110011010011001100110010110011011001100110011001100110011001100,
64'b0011001100110011110011001100110001011010010110100101101001011010,
64'b1111111100000000111111110000000011001100001100110011001111001100,
64'b0101101010100101101001010101101000001111000011111111000011110000,
64'b1001100101100110100110010110011001101001011010011001011010010110,
64'b1001011010010110100101101001011010101010101010101010101010101010,
64'b1001011001101001011010011001011000001111000011111111000011110000,
64'b0101010110101010010101011010101000001111111100000000111111110000,
64'b0110011001100110011001100110011011110000111100001111000011110000,
64'b1001011001101001011010011001011001100110100110011001100101100110,
64'b1100001100111100110000110011110010011001011001101001100101100110,
64'b1001011001101001011010011001011011111111111111110000000000000000,
64'b0000000011111111111111110000000000001111000011111111000011110000,
64'b1010101001010101010101011010101011110000111100001111000011110000,
64'b0101101010100101101001010101101000110011110011000011001111001100,
64'b0110011010011001100110010110011000001111000011111111000011110000,
64'b1001100110011001011001100110011001010101101010100101010110101010,
64'b1001100101100110100110010110011001101001100101100110100110010110,
64'b1010010101011010101001010101101001100110011001100110011001100110,
64'b0000111100001111111100001111000011111111000000001111111100000000,
64'b0000000011111111111111110000000010101010010101010101010110101010,
64'b1001011001101001011010011001011011111111000000001111111100000000,
64'b0000000000000000000000000000000011000011110000110011110000111100,
64'b1111000011110000111100001111000001101001011010011001011010010110,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1100001111000011001111000011110001010101101010100101010110101010,
64'b1111000000001111000011111111000001010101101010100101010110101010,
64'b0110011001100110011001100110011000001111000011111111000011110000,
64'b0101101010100101101001010101101011111111000000001111111100000000,
64'b1100001100111100110000110011110010011001100110010110011001100110,
64'b1001100101100110100110010110011000111100110000111100001100111100,
64'b0101010110101010010101011010101000111100001111000011110000111100,
64'b1111111100000000111111110000000011001100001100110011001111001100,
64'b0101010101010101101010101010101010101010010101010101010110101010,
64'b1001011001101001011010011001011011111111000000001111111100000000,
64'b1010101010101010101010101010101000110011001100111100110011001100,
64'b1111111100000000111111110000000011000011110000110011110000111100,
64'b0000000000000000000000000000000010010110011010010110100110010110,
64'b0000111111110000000011111111000010100101101001010101101001011010,
64'b1010101001010101010101011010101001011010101001011010010101011010,
64'b1001011010010110100101101001011011111111111111110000000000000000,
64'b1100110000110011001100111100110001100110100110011001100101100110,
64'b0101101010100101101001010101101001101001100101100110100110010110,
64'b1100001111000011001111000011110010101010101010101010101010101010,
64'b1100110011001100110011001100110011000011001111001100001100111100,
64'b0110011010011001100110010110011010010110011010010110100110010110,
64'b0101010110101010010101011010101000000000111111111111111100000000,
64'b0011110000111100001111000011110011111111000000001111111100000000,
64'b0101101010100101101001010101101011001100001100110011001111001100,
64'b0101010110101010010101011010101000001111000011111111000011110000,
64'b0011110011000011110000110011110010101010101010101010101010101010,
64'b1001011001101001011010011001011000001111111100000000111111110000,
64'b0101101010100101101001010101101000001111000011111111000011110000,
64'b0110100101101001100101101001011010101010010101010101010110101010,
64'b0011110011000011110000110011110001011010101001011010010101011010,
64'b0011001100110011110011001100110011000011110000110011110000111100,
64'b0101010101010101101010101010101000111100110000111100001100111100,
64'b0011110000111100001111000011110001101001100101100110100110010110,
64'b0101101010100101101001010101101010010110011010010110100110010110,
64'b0000000011111111111111110000000001010101010101011010101010101010,
64'b1010010110100101010110100101101001010101010101011010101010101010,
64'b1111000011110000111100001111000000001111000011111111000011110000,
64'b0011001111001100001100111100110001010101101010100101010110101010,
64'b1100110011001100110011001100110001100110011001100110011001100110,
64'b0000000011111111111111110000000000000000111111111111111100000000,
64'b0000111100001111111100001111000011111111000000001111111100000000,
64'b0110100101101001100101101001011010011001100110010110011001100110,
64'b0110100101101001100101101001011001100110100110011001100101100110,
64'b0000111111110000000011111111000010100101010110101010010101011010,
64'b1001011001101001011010011001011001011010101001011010010101011010,
64'b1100001100111100110000110011110001101001100101100110100110010110,
64'b1100110000110011001100111100110010010110011010010110100110010110,
64'b0101010101010101101010101010101001100110011001100110011001100110,
64'b1001100101100110100110010110011001100110011001100110011001100110,
64'b0101010110101010010101011010101001010101101010100101010110101010,
64'b0000111100001111111100001111000010011001100110010110011001100110,
64'b1111000011110000111100001111000000111100001111000011110000111100,
64'b1111111111111111000000000000000011111111111111110000000000000000,
64'b0101010110101010010101011010101001010101010101011010101010101010,
64'b0110100110010110011010011001011000111100001111000011110000111100,
64'b0110100110010110011010011001011001101001011010011001011010010110,
64'b1010101001010101010101011010101001100110100110011001100101100110,
64'b0011110011000011110000110011110011001100001100110011001111001100,
64'b1010010101011010101001010101101001101001100101100110100110010110,
64'b0011110011000011110000110011110010100101101001010101101001011010,
64'b1111111100000000111111110000000000001111111100000000111111110000,
64'b1100001100111100110000110011110010010110011010010110100110010110,
64'b0000111111110000000011111111000000001111111100000000111111110000,
64'b0101010101010101101010101010101010010110011010010110100110010110,
64'b0110100101101001100101101001011010011001100110010110011001100110,
64'b1001011010010110100101101001011010010110100101101001011010010110,
64'b1111000000001111000011111111000000001111111100000000111111110000,
64'b0011110000111100001111000011110010100101101001010101101001011010,
64'b0000111100001111111100001111000011110000111100001111000011110000,
64'b0110011010011001100110010110011000111100110000111100001100111100,
64'b1010101010101010101010101010101001010101101010100101010110101010,
64'b1111111100000000111111110000000000001111111100000000111111110000,
64'b1100001111000011001111000011110010011001011001101001100101100110,
64'b1100110000110011001100111100110010101010010101010101010110101010,
64'b0101101001011010010110100101101000111100110000111100001100111100,
64'b0011110000111100001111000011110010101010010101010101010110101010,
64'b0110011010011001100110010110011000111100110000111100001100111100,
64'b0101010101010101101010101010101010010110100101101001011010010110,
64'b1111111100000000111111110000000001101001100101100110100110010110,
64'b0110100101101001100101101001011000000000111111111111111100000000,
64'b1010010110100101010110100101101000110011110011000011001111001100,
64'b1100110011001100110011001100110001010101101010100101010110101010,
64'b0011110011000011110000110011110011110000000011110000111111110000,
64'b1001011001101001011010011001011010011001100110010110011001100110,
64'b0110011001100110011001100110011011111111000000001111111100000000,
64'b1001011010010110100101101001011011000011110000110011110000111100,
64'b0011110011000011110000110011110000110011001100111100110011001100,
64'b0011001100110011110011001100110001011010101001011010010101011010,
64'b0011001100110011110011001100110010011001100110010110011001100110,
64'b0110100110010110011010011001011001011010101001011010010101011010,
64'b0101101010100101101001010101101001101001100101100110100110010110,
64'b1100001111000011001111000011110000111100110000111100001100111100,
64'b1010101010101010101010101010101011111111111111110000000000000000,
64'b1001100110011001011001100110011010100101101001010101101001011010,
64'b0110100110010110011010011001011000110011001100111100110011001100,
64'b1010010110100101010110100101101000000000111111111111111100000000,
64'b0110011001100110011001100110011010010110100101101001011010010110,
64'b1111000011110000111100001111000010101010101010101010101010101010,
64'b1100001100111100110000110011110010100101010110101010010101011010,
64'b1111000000001111000011111111000001011010010110100101101001011010,
64'b0101101001011010010110100101101001100110100110011001100101100110,
64'b0101101001011010010110100101101010010110100101101001011010010110,
64'b1001011001101001011010011001011001100110100110011001100101100110,
64'b1100110000110011001100111100110010010110011010010110100110010110,
64'b1010010101011010101001010101101011110000000011110000111111110000,
64'b0110011001100110011001100110011010101010101010101010101010101010,
64'b0011110000111100001111000011110010011001011001101001100101100110,
64'b1001011001101001011010011001011001011010010110100101101001011010,
64'b0011001111001100001100111100110001010101010101011010101010101010,
64'b1001011010010110100101101001011001101001100101100110100110010110,
64'b1111111100000000111111110000000011001100110011001100110011001100,
64'b1111000000001111000011111111000011001100001100110011001111001100,
64'b0000000011111111111111110000000000110011110011000011001111001100,
64'b1001100101100110100110010110011011000011110000110011110000111100,
64'b0011001111001100001100111100110001101001100101100110100110010110,
64'b0011110011000011110000110011110011000011110000110011110000111100,
64'b1010010110100101010110100101101010010110011010010110100110010110,
64'b0110011010011001100110010110011010101010010101010101010110101010,
64'b0011110000111100001111000011110001100110011001100110011001100110,
64'b0000111111110000000011111111000011000011110000110011110000111100,
64'b0011110011000011110000110011110000110011110011000011001111001100,
64'b1010010110100101010110100101101011001100110011001100110011001100,
64'b1100001100111100110000110011110010010110011010010110100110010110,
64'b0000000000000000000000000000000011110000111100001111000011110000,
64'b1010101001010101010101011010101010100101101001010101101001011010,
64'b0101010101010101101010101010101010100101101001010101101001011010,
64'b0110100101101001100101101001011000001111111100000000111111110000,
64'b0000111100001111111100001111000010010110011010010110100110010110,
64'b1111000000001111000011111111000000001111111100000000111111110000,
64'b1001100101100110100110010110011010010110011010010110100110010110,
64'b0110100101101001100101101001011010011001100110010110011001100110,
64'b1010010101011010101001010101101010010110100101101001011010010110,
64'b0000000011111111111111110000000000001111111100000000111111110000,
64'b1111000000001111000011111111000010100101101001010101101001011010,
64'b1001100101100110100110010110011011110000111100001111000011110000,
64'b0101101010100101101001010101101000111100110000111100001100111100,
64'b0000000000000000000000000000000001010101101010100101010110101010,
64'b0101010101010101101010101010101001011010010110100101101001011010,
64'b1010010101011010101001010101101010101010010101010101010110101010,
64'b1100110000110011001100111100110001100110011001100110011001100110,
64'b1010010110100101010110100101101010100101101001010101101001011010,
64'b0011110011000011110000110011110000001111000011111111000011110000,
64'b0101101001011010010110100101101001010101101010100101010110101010,
64'b0000000000000000000000000000000001101001100101100110100110010110,
64'b1100001100111100110000110011110010100101010110101010010101011010,
64'b0110100110010110011010011001011011000011110000110011110000111100,
64'b1010101001010101010101011010101001101001011010011001011010010110,
64'b1111111111111111000000000000000010100101010110101010010101011010,
64'b0000000011111111111111110000000011001100001100110011001111001100,
64'b0011110000111100001111000011110000110011110011000011001111001100,
64'b1001100110011001011001100110011000110011110011000011001111001100,
64'b1100001111000011001111000011110000110011001100111100110011001100,
64'b1100001100111100110000110011110010010110100101101001011010010110,
64'b0011110011000011110000110011110000110011110011000011001111001100,
64'b0110011001100110011001100110011001010101101010100101010110101010,
64'b1100001100111100110000110011110010011001100110010110011001100110,
64'b0000000000000000000000000000000000111100110000111100001100111100,
64'b0011001100110011110011001100110011001100001100110011001111001100,
64'b0101010101010101101010101010101000001111111100000000111111110000,
64'b1001100101100110100110010110011001101001100101100110100110010110,
64'b0101010101010101101010101010101001100110100110011001100101100110,
64'b0101010110101010010101011010101000001111000011111111000011110000,
64'b1001100101100110100110010110011001011010010110100101101001011010,
64'b0110100101101001100101101001011000001111000011111111000011110000,
64'b0000000000000000000000000000000011110000111100001111000011110000,
64'b1001011010010110100101101001011001101001100101100110100110010110,
64'b0101010110101010010101011010101000001111000011111111000011110000,
64'b1010101001010101010101011010101000110011001100111100110011001100,
64'b1010101001010101010101011010101000111100001111000011110000111100,
64'b0000000000000000000000000000000001011010101001011010010101011010,
64'b0011001111001100001100111100110010100101101001010101101001011010,
64'b0000111111110000000011111111000010101010010101010101010110101010,
64'b1100001100111100110000110011110000111100110000111100001100111100,
64'b0011001100110011110011001100110011000011110000110011110000111100,
64'b1001100101100110100110010110011001010101101010100101010110101010,
64'b0000000000000000000000000000000010011001011001101001100101100110,
64'b0110100110010110011010011001011001010101101010100101010110101010,
64'b1010101010101010101010101010101001010101101010100101010110101010,
64'b1100001100111100110000110011110000111100110000111100001100111100,
64'b0011001100110011110011001100110011111111000000001111111100000000,
64'b0011001100110011110011001100110001011010010110100101101001011010,
64'b1001100110011001011001100110011010100101010110101010010101011010,
64'b1010101010101010101010101010101011001100001100110011001111001100,
64'b0000111100001111111100001111000010011001011001101001100101100110,
64'b0000000011111111111111110000000010011001100110010110011001100110,
64'b1111000000001111000011111111000001011010101001011010010101011010,
64'b1111000011110000111100001111000010100101010110101010010101011010,
64'b0110100101101001100101101001011010011001100110010110011001100110,
64'b0000000000000000000000000000000000111100001111000011110000111100,
64'b0110100110010110011010011001011000110011001100111100110011001100,
64'b0110100110010110011010011001011000110011001100111100110011001100,
64'b0011110000111100001111000011110011110000000011110000111111110000,
64'b0101010101010101101010101010101001010101010101011010101010101010,
64'b0110011010011001100110010110011000110011110011000011001111001100,
64'b1100110011001100110011001100110011001100001100110011001111001100,
64'b0110011001100110011001100110011000001111000011111111000011110000,
64'b0011110000111100001111000011110001101001011010011001011010010110,
64'b0011110011000011110000110011110000111100001111000011110000111100,
64'b0000000000000000000000000000000001100110100110011001100101100110,
64'b1010101001010101010101011010101001100110100110011001100101100110,
64'b1100001111000011001111000011110000111100001111000011110000111100,
64'b1001011010010110100101101001011010100101010110101010010101011010,
64'b1100001100111100110000110011110011110000111100001111000011110000,
64'b1001100110011001011001100110011001011010010110100101101001011010,
64'b1100001111000011001111000011110010101010010101010101010110101010,
64'b0110100101101001100101101001011001100110011001100110011001100110,
64'b0101010110101010010101011010101010100101101001010101101001011010,
64'b0000000000000000000000000000000000001111000011111111000011110000,
64'b0011110000111100001111000011110001010101101010100101010110101010,
64'b1100110011001100110011001100110001101001100101100110100110010110,
64'b1001100110011001011001100110011010100101010110101010010101011010,
64'b0000000011111111111111110000000011000011110000110011110000111100,
64'b1100110011001100110011001100110001101001011010011001011010010110,
64'b1010010110100101010110100101101010100101010110101010010101011010,
64'b0101010110101010010101011010101000110011110011000011001111001100,
64'b0101101010100101101001010101101010101010010101010101010110101010,
64'b0011110000111100001111000011110010010110100101101001011010010110,
64'b1010010101011010101001010101101011111111000000001111111100000000,
64'b0110100110010110011010011001011000110011001100111100110011001100,
64'b1001100110011001011001100110011000001111000011111111000011110000,
64'b0000000000000000000000000000000000001111111100000000111111110000,
64'b0000111111110000000011111111000010011001100110010110011001100110,
64'b1111000011110000111100001111000011111111111111110000000000000000,
64'b0011110000111100001111000011110010100101101001010101101001011010,
64'b0101010101010101101010101010101010100101101001010101101001011010,
64'b0101101001011010010110100101101010010110011010010110100110010110,
64'b0011001111001100001100111100110001100110011001100110011001100110,
64'b0110011001100110011001100110011011001100110011001100110011001100,
64'b1001100101100110100110010110011011001100110011001100110011001100,
64'b0000000000000000000000000000000011001100110011001100110011001100,
64'b0000000000000000000000000000000000110011110011000011001111001100,
64'b1001100101100110100110010110011001010101010101011010101010101010,
64'b0000000011111111111111110000000001101001011010011001011010010110,
64'b1111000011110000111100001111000011110000000011110000111111110000,
64'b0000000011111111111111110000000000111100001111000011110000111100,
64'b0011110000111100001111000011110001101001100101100110100110010110,
64'b0110011001100110011001100110011011110000111100001111000011110000,
64'b0110011010011001100110010110011000110011001100111100110011001100,
64'b0110011010011001100110010110011001101001100101100110100110010110,
64'b0000111111110000000011111111000010010110011010010110100110010110,
64'b0000000000000000000000000000000011001100110011001100110011001100,
64'b1001011010010110100101101001011001011010010110100101101001011010,
64'b1010010101011010101001010101101011110000111100001111000011110000,
64'b1100110000110011001100111100110000001111000011111111000011110000,
64'b0110011001100110011001100110011011001100110011001100110011001100,
64'b1100001100111100110000110011110001101001100101100110100110010110,
64'b0000111111110000000011111111000010101010010101010101010110101010,
64'b1111111111111111000000000000000010100101010110101010010101011010,
64'b0110011001100110011001100110011000111100110000111100001100111100,
64'b0101010110101010010101011010101011111111000000001111111100000000,
64'b0110100110010110011010011001011011110000111100001111000011110000,
64'b1001011010010110100101101001011010010110011010010110100110010110,
64'b1010101010101010101010101010101000111100110000111100001100111100,
64'b0011110000111100001111000011110001011010010110100101101001011010,
64'b0110100110010110011010011001011010011001011001101001100101100110,
64'b1100110000110011001100111100110011111111000000001111111100000000,
64'b0000111100001111111100001111000011111111000000001111111100000000,
64'b1001011010010110100101101001011001011010010110100101101001011010,
64'b1111000000001111000011111111000000111100110000111100001100111100,
64'b0000000011111111111111110000000000110011001100111100110011001100,
64'b0000000000000000000000000000000001100110100110011001100101100110,
64'b1001011010010110100101101001011011110000000011110000111111110000,
64'b0011001100110011110011001100110001010101010101011010101010101010,
64'b0011110011000011110000110011110011111111000000001111111100000000,
64'b1100001100111100110000110011110000111100110000111100001100111100,
64'b1100110011001100110011001100110001011010101001011010010101011010,
64'b0000111111110000000011111111000010011001011001101001100101100110,
64'b1100001100111100110000110011110000111100001111000011110000111100,
64'b1010101001010101010101011010101001011010101001011010010101011010,
64'b1001100110011001011001100110011000110011110011000011001111001100,
64'b1100110000110011001100111100110010010110011010010110100110010110,
64'b0011110000111100001111000011110011001100110011001100110011001100,
64'b0000111100001111111100001111000000000000000000000000000000000000,
64'b1010101010101010101010101010101001101001011010011001011010010110,
64'b0000000000000000000000000000000001101001011010011001011010010110,
64'b1001100101100110100110010110011000001111111100000000111111110000,
64'b1111000011110000111100001111000011111111000000001111111100000000,
64'b1010010101011010101001010101101000001111111100000000111111110000,
64'b1111000000001111000011111111000001100110011001100110011001100110,
64'b1100001100111100110000110011110010101010101010101010101010101010,
64'b0000111111110000000011111111000010100101010110101010010101011010,
64'b1001011001101001011010011001011011001100001100110011001111001100,
64'b0101101010100101101001010101101010100101101001010101101001011010,
64'b0000000000000000000000000000000000111100110000111100001100111100,
64'b1001100110011001011001100110011001011010010110100101101001011010,
64'b1010010101011010101001010101101000000000000000000000000000000000,
64'b0110011001100110011001100110011011000011001111001100001100111100,
64'b1100001100111100110000110011110001101001100101100110100110010110,
64'b1010101001010101010101011010101010101010010101010101010110101010,
64'b0101010101010101101010101010101011111111111111110000000000000000,
64'b0011001111001100001100111100110000000000111111111111111100000000,
64'b0000000000000000000000000000000000111100001111000011110000111100,
64'b1001100101100110100110010110011011001100110011001100110011001100,
64'b0101010110101010010101011010101001100110100110011001100101100110,
64'b1001100110011001011001100110011000001111000011111111000011110000,
64'b1010101010101010101010101010101010011001011001101001100101100110,
64'b0000111100001111111100001111000001011010101001011010010101011010,
64'b0000000011111111111111110000000010011001011001101001100101100110,
64'b0011110011000011110000110011110000000000000000000000000000000000,
64'b0011110000111100001111000011110011110000000011110000111111110000,
64'b0011001100110011110011001100110000111100110000111100001100111100,
64'b0101101010100101101001010101101000110011001100111100110011001100,
64'b1100110000110011001100111100110010101010101010101010101010101010,
64'b0101101001011010010110100101101001010101010101011010101010101010,
64'b0000000011111111111111110000000010100101010110101010010101011010,
64'b0000000000000000000000000000000011110000111100001111000011110000,
64'b0011001100110011110011001100110011000011110000110011110000111100,
64'b0011110000111100001111000011110001010101101010100101010110101010,
64'b0110011001100110011001100110011001101001011010011001011010010110,
64'b1111111100000000111111110000000011001100001100110011001111001100,
64'b0101010101010101101010101010101001101001011010011001011010010110,
64'b0101101010100101101001010101101000000000000000000000000000000000,
64'b1010010101011010101001010101101000000000111111111111111100000000,
64'b1111000011110000111100001111000001011010101001011010010101011010,
64'b0110011010011001100110010110011001011010010110100101101001011010,
64'b1010010110100101010110100101101001100110011001100110011001100110,
64'b1001100101100110100110010110011011001100110011001100110011001100,
64'b1111111111111111000000000000000001100110100110011001100101100110,
64'b1010101010101010101010101010101011111111000000001111111100000000,
64'b0101101001011010010110100101101000001111111100000000111111110000,
64'b1010010101011010101001010101101010011001100110010110011001100110,
64'b0011110000111100001111000011110011000011001111001100001100111100,
64'b1111111111111111000000000000000010100101101001010101101001011010,
64'b1100110011001100110011001100110001101001100101100110100110010110,
64'b0110011010011001100110010110011010101010101010101010101010101010,
64'b0110011010011001100110010110011011111111111111110000000000000000,
64'b1111111100000000111111110000000001100110100110011001100101100110,
64'b1100001111000011001111000011110010011001011001101001100101100110,
64'b1001100101100110100110010110011000111100001111000011110000111100,
64'b0110100101101001100101101001011011110000111100001111000011110000,
64'b0000000000000000000000000000000011000011110000110011110000111100,
64'b0110011001100110011001100110011010101010101010101010101010101010,
64'b0011001111001100001100111100110000000000111111111111111100000000,
64'b1100110000110011001100111100110000111100001111000011110000111100,
64'b0000111111110000000011111111000001011010101001011010010101011010,
64'b0000000000000000000000000000000000110011110011000011001111001100,
64'b0101101001011010010110100101101010010110011010010110100110010110,
64'b1100001111000011001111000011110011001100110011001100110011001100,
64'b0110100101101001100101101001011000000000000000000000000000000000,
64'b0101010101010101101010101010101001101001011010011001011010010110,
64'b0000111111110000000011111111000001101001011010011001011010010110,
64'b0110100101101001100101101001011000001111111100000000111111110000,
64'b1100001100111100110000110011110011111111000000001111111100000000,
64'b1010101010101010101010101010101000001111111100000000111111110000,
64'b0011110000111100001111000011110001100110011001100110011001100110,
64'b1111000011110000111100001111000000001111000011111111000011110000,
64'b0011001111001100001100111100110010010110100101101001011010010110,
64'b1010101001010101010101011010101011111111000000001111111100000000,
64'b1111000011110000111100001111000011000011001111001100001100111100,
64'b1001100110011001011001100110011011001100001100110011001111001100,
64'b0000000000000000000000000000000000110011110011000011001111001100,
64'b1001011010010110100101101001011011000011001111001100001100111100,
64'b0011001111001100001100111100110001101001011010011001011010010110,
64'b0101101001011010010110100101101010010110011010010110100110010110,
64'b0101010110101010010101011010101001011010101001011010010101011010,
64'b1001100101100110100110010110011010011001011001101001100101100110,
64'b0000111100001111111100001111000001010101101010100101010110101010,
64'b1010010101011010101001010101101011111111000000001111111100000000,
64'b0000111111110000000011111111000001010101101010100101010110101010,
64'b0011110011000011110000110011110001101001100101100110100110010110,
64'b1001100101100110100110010110011011111111111111110000000000000000,
64'b1010010101011010101001010101101011110000000011110000111111110000,
64'b1010010110100101010110100101101000001111000011111111000011110000,
64'b1010101010101010101010101010101010100101101001010101101001011010,
64'b0101010110101010010101011010101011110000000011110000111111110000,
64'b0011110011000011110000110011110011000011001111001100001100111100,
64'b0110100110010110011010011001011010010110011010010110100110010110,
64'b0110011010011001100110010110011001100110100110011001100101100110,
64'b0101101010100101101001010101101001101001011010011001011010010110,
64'b1111000000001111000011111111000000110011001100111100110011001100,
64'b0011110000111100001111000011110000000000000000000000000000000000,
64'b0101101010100101101001010101101000110011001100111100110011001100,
64'b1100001111000011001111000011110000111100110000111100001100111100,
64'b1100001100111100110000110011110000000000000000000000000000000000,
64'b0011110011000011110000110011110010101010010101010101010110101010,
64'b1010101001010101010101011010101001010101101010100101010110101010,
64'b0110011001100110011001100110011010011001011001101001100101100110,
64'b1010010110100101010110100101101010101010010101010101010110101010,
64'b1100001111000011001111000011110001011010101001011010010101011010,
64'b1100110000110011001100111100110000111100110000111100001100111100,
64'b1001011001101001011010011001011001101001011010011001011010010110,
64'b1111111111111111000000000000000001101001100101100110100110010110,
64'b1010010101011010101001010101101001011010010110100101101001011010,
64'b0000000000000000000000000000000010101010101010101010101010101010,
64'b1100110000110011001100111100110001011010010110100101101001011010,
64'b1010010101011010101001010101101001011010101001011010010101011010,
64'b0101101010100101101001010101101010101010101010101010101010101010,
64'b1111000000001111000011111111000000110011001100111100110011001100,
64'b1001100110011001011001100110011010011001100110010110011001100110,
64'b1001011010010110100101101001011011000011110000110011110000111100,
64'b0011001111001100001100111100110000110011001100111100110011001100,
64'b1010010101011010101001010101101001100110100110011001100101100110,
64'b1010010110100101010110100101101001011010101001011010010101011010,
64'b1001011001101001011010011001011001101001100101100110100110010110,
64'b1010101010101010101010101010101010010110011010010110100110010110,
64'b0110011010011001100110010110011000110011110011000011001111001100,
64'b0000000000000000000000000000000011001100110011001100110011001100,
64'b1111111111111111000000000000000000110011110011000011001111001100,
64'b0101010101010101101010101010101011001100001100110011001111001100,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b0101101010100101101001010101101011110000111100001111000011110000,
64'b0000111100001111111100001111000010010110100101101001011010010110,
64'b0110100110010110011010011001011010100101010110101010010101011010,
64'b1001100110011001011001100110011001011010010110100101101001011010,
64'b1111111111111111000000000000000001101001011010011001011010010110,
64'b0110100110010110011010011001011001100110100110011001100101100110,
64'b1100001111000011001111000011110010010110011010010110100110010110,
64'b1111111100000000111111110000000000111100110000111100001100111100,
64'b1100110011001100110011001100110010100101101001010101101001011010,
64'b0000111111110000000011111111000011110000111100001111000011110000,
64'b1111000011110000111100001111000010100101101001010101101001011010,
64'b0101010110101010010101011010101000001111000011111111000011110000,
64'b0011110011000011110000110011110010010110100101101001011010010110,
64'b0011110011000011110000110011110011111111000000001111111100000000,
64'b1100110000110011001100111100110011000011001111001100001100111100,
64'b1001011001101001011010011001011011001100001100110011001111001100,
64'b1010101010101010101010101010101000110011110011000011001111001100,
64'b1001100101100110100110010110011011000011001111001100001100111100,
64'b1100110000110011001100111100110001101001011010011001011010010110,
64'b0101101001011010010110100101101010010110011010010110100110010110,
64'b1100110000110011001100111100110001011010101001011010010101011010,
64'b1111111111111111000000000000000010011001011001101001100101100110,
64'b0101101001011010010110100101101001010101101010100101010110101010,
64'b0101010110101010010101011010101001101001100101100110100110010110,
64'b0011001100110011110011001100110001100110011001100110011001100110,
64'b1111000000001111000011111111000011000011110000110011110000111100,
64'b0101101010100101101001010101101000001111000011111111000011110000,
64'b1010010110100101010110100101101001101001100101100110100110010110,
64'b1001011001101001011010011001011000001111000011111111000011110000,
64'b0110011001100110011001100110011000110011001100111100110011001100,
64'b1100001111000011001111000011110011000011110000110011110000111100,
64'b0000111100001111111100001111000010011001011001101001100101100110,
64'b1001100101100110100110010110011011000011110000110011110000111100,
64'b0000111100001111111100001111000011111111111111110000000000000000,
64'b1010101010101010101010101010101001100110011001100110011001100110,
64'b1001100101100110100110010110011001101001100101100110100110010110,
64'b1100001111000011001111000011110011001100001100110011001111001100,
64'b1100001100111100110000110011110000001111111100000000111111110000,
64'b0000000000000000000000000000000010100101101001010101101001011010,
64'b1001011001101001011010011001011010100101010110101010010101011010,
64'b0000000011111111111111110000000000001111111100000000111111110000,
64'b1001011001101001011010011001011011111111000000001111111100000000,
64'b0000000000000000000000000000000011001100110011001100110011001100,
64'b0011110000111100001111000011110010010110100101101001011010010110,
64'b0000111111110000000011111111000000110011001100111100110011001100,
64'b0011110011000011110000110011110001011010010110100101101001011010,
64'b0110011001100110011001100110011000110011110011000011001111001100,
64'b0110100101101001100101101001011010011001100110010110011001100110,
64'b1001100101100110100110010110011001100110011001100110011001100110,
64'b1111111100000000111111110000000000001111000011111111000011110000,
64'b0110100101101001100101101001011010101010010101010101010110101010,
64'b1010101001010101010101011010101000110011110011000011001111001100,
64'b1100110000110011001100111100110001100110100110011001100101100110,
64'b1100110011001100110011001100110000000000111111111111111100000000,
64'b1001011001101001011010011001011011111111111111110000000000000000,
64'b0011110000111100001111000011110011110000111100001111000011110000,
64'b0011110000111100001111000011110011000011001111001100001100111100,
64'b0101101010100101101001010101101011110000111100001111000011110000,
64'b1010010110100101010110100101101010011001011001101001100101100110,
64'b0000111111110000000011111111000000001111000011111111000011110000,
64'b1100110000110011001100111100110000111100001111000011110000111100,
64'b0011001111001100001100111100110010010110100101101001011010010110,
64'b1111111111111111000000000000000011111111000000001111111100000000,
64'b1100001100111100110000110011110010011001100110010110011001100110,
64'b1001100110011001011001100110011010100101101001010101101001011010,
64'b1010010110100101010110100101101011000011110000110011110000111100,
64'b0101101001011010010110100101101001010101010101011010101010101010,
64'b0011110011000011110000110011110010101010101010101010101010101010,
64'b1010010101011010101001010101101001010101101010100101010110101010,
64'b0000111111110000000011111111000011110000000011110000111111110000,
64'b1100110000110011001100111100110011111111000000001111111100000000,
64'b1001100101100110100110010110011011000011110000110011110000111100,
64'b1010101001010101010101011010101011111111000000001111111100000000,
64'b0000111100001111111100001111000010100101010110101010010101011010,
64'b0101101001011010010110100101101011000011001111001100001100111100,
64'b0101101001011010010110100101101010100101101001010101101001011010,
64'b0110100101101001100101101001011000001111111100000000111111110000,
64'b1001011001101001011010011001011000110011001100111100110011001100,
64'b0110100110010110011010011001011001010101101010100101010110101010,
64'b0000000011111111111111110000000011111111111111110000000000000000,
64'b1111000000001111000011111111000001100110011001100110011001100110,
64'b1111000000001111000011111111000010100101101001010101101001011010,
64'b0011001100110011110011001100110000110011001100111100110011001100,
64'b0101010101010101101010101010101000001111000011111111000011110000,
64'b0011110011000011110000110011110001011010010110100101101001011010,
64'b1010101001010101010101011010101011001100001100110011001111001100,
64'b0101101010100101101001010101101011000011001111001100001100111100,
64'b0011110000111100001111000011110010101010101010101010101010101010,
64'b0110100110010110011010011001011000110011110011000011001111001100,
64'b1111000011110000111100001111000010101010010101010101010110101010,
64'b0011110000111100001111000011110011110000111100001111000011110000,
64'b0110011010011001100110010110011010011001100110010110011001100110,
64'b0110011001100110011001100110011000000000000000000000000000000000,
64'b1010101001010101010101011010101010010110100101101001011010010110,
64'b0011110011000011110000110011110000110011110011000011001111001100,
64'b0110100110010110011010011001011001011010010110100101101001011010,
64'b0011110000111100001111000011110001010101101010100101010110101010,
64'b0000111100001111111100001111000010011001011001101001100101100110,
64'b0000000011111111111111110000000000001111000011111111000011110000,
64'b0110100110010110011010011001011001011010101001011010010101011010,
64'b0000000000000000000000000000000011001100110011001100110011001100,
64'b0110011010011001100110010110011000001111000011111111000011110000,
64'b1100110011001100110011001100110000110011001100111100110011001100,
64'b1010010110100101010110100101101001010101101010100101010110101010,
64'b0011001100110011110011001100110000111100001111000011110000111100,
64'b0000111100001111111100001111000010101010101010101010101010101010,
64'b0011001100110011110011001100110011000011001111001100001100111100,
64'b1100110000110011001100111100110000001111000011111111000011110000,
64'b1010010110100101010110100101101000110011110011000011001111001100,
64'b0101010110101010010101011010101000110011001100111100110011001100,
64'b1010101010101010101010101010101011000011110000110011110000111100,
64'b1100110000110011001100111100110011111111000000001111111100000000,
64'b1001100101100110100110010110011001100110100110011001100101100110,
64'b1010010101011010101001010101101001011010010110100101101001011010,
64'b1100001111000011001111000011110011111111000000001111111100000000,
64'b0101101001011010010110100101101001011010010110100101101001011010,
64'b0011001111001100001100111100110010011001100110010110011001100110,
64'b0101101001011010010110100101101000001111111100000000111111110000,
64'b0101010110101010010101011010101011001100110011001100110011001100,
64'b0101101001011010010110100101101011110000000011110000111111110000,
64'b1010010110100101010110100101101011111111000000001111111100000000,
64'b1001100101100110100110010110011010100101101001010101101001011010,
64'b1001100110011001011001100110011011110000111100001111000011110000,
64'b1100110011001100110011001100110010100101010110101010010101011010,
64'b0000111100001111111100001111000001010101010101011010101010101010,
64'b0110100101101001100101101001011011000011110000110011110000111100,
64'b0011001111001100001100111100110010011001011001101001100101100110,
64'b0000111111110000000011111111000001010101010101011010101010101010,
64'b1001100101100110100110010110011000110011110011000011001111001100,
64'b0000111100001111111100001111000000111100001111000011110000111100,
64'b0011001111001100001100111100110010101010010101010101010110101010,
64'b0011001100110011110011001100110011110000111100001111000011110000,
64'b0011001111001100001100111100110000000000111111111111111100000000,
64'b0011001111001100001100111100110001010101010101011010101010101010,
64'b0110100101101001100101101001011000110011110011000011001111001100,
64'b0011110000111100001111000011110001010101101010100101010110101010,
64'b0101101001011010010110100101101011001100001100110011001111001100,
64'b1111111100000000111111110000000011001100110011001100110011001100,
64'b0110100110010110011010011001011010100101010110101010010101011010,
64'b0101101001011010010110100101101010010110100101101001011010010110,
64'b0000000011111111111111110000000011001100110011001100110011001100,
64'b1100001111000011001111000011110010100101101001010101101001011010,
64'b1111111100000000111111110000000000001111111100000000111111110000,
64'b1010010110100101010110100101101000110011001100111100110011001100,
64'b1111000011110000111100001111000001010101101010100101010110101010,
64'b1010010110100101010110100101101011111111111111110000000000000000,
64'b0000111100001111111100001111000001100110011001100110011001100110,
64'b1100001100111100110000110011110010100101101001010101101001011010,
64'b1010010101011010101001010101101000110011001100111100110011001100,
64'b0011001111001100001100111100110000001111000011111111000011110000,
64'b1111111111111111000000000000000001011010010110100101101001011010,
64'b0011110011000011110000110011110011001100001100110011001111001100,
64'b0011001111001100001100111100110011000011001111001100001100111100,
64'b0101101001011010010110100101101000000000111111111111111100000000,
64'b1111111100000000111111110000000010101010101010101010101010101010,
64'b1100001111000011001111000011110001011010010110100101101001011010,
64'b0101010101010101101010101010101011001100001100110011001111001100,
64'b1010010101011010101001010101101000000000111111111111111100000000,
64'b0000000011111111111111110000000000000000111111111111111100000000,
64'b0110100110010110011010011001011010101010010101010101010110101010,
64'b0011001111001100001100111100110000111100110000111100001100111100,
64'b1010010101011010101001010101101000111100001111000011110000111100,
64'b1100001111000011001111000011110000110011001100111100110011001100,
64'b1100110000110011001100111100110011001100001100110011001111001100,
64'b0101101001011010010110100101101010100101010110101010010101011010,
64'b1111111100000000111111110000000001010101101010100101010110101010,
64'b1100001100111100110000110011110001010101010101011010101010101010,
64'b0000000011111111111111110000000001100110011001100110011001100110,
64'b1100110000110011001100111100110000110011110011000011001111001100,
64'b0011001100110011110011001100110000001111000011111111000011110000,
64'b1100001111000011001111000011110001010101010101011010101010101010,
64'b1111111100000000111111110000000001010101010101011010101010101010,
64'b1111111111111111000000000000000010011001100110010110011001100110,
64'b0011110011000011110000110011110001011010101001011010010101011010,
64'b0110100101101001100101101001011010100101010110101010010101011010,
64'b1100110000110011001100111100110011110000111100001111000011110000,
64'b0110100110010110011010011001011010100101101001010101101001011010,
64'b1100001100111100110000110011110001100110100110011001100101100110,
64'b1111111100000000111111110000000011001100110011001100110011001100,
64'b1010101001010101010101011010101011001100110011001100110011001100,
64'b0000000011111111111111110000000010010110100101101001011010010110,
64'b0110011001100110011001100110011000001111000011111111000011110000,
64'b0000111100001111111100001111000011111111000000001111111100000000,
64'b0000000000000000000000000000000001100110011001100110011001100110,
64'b0101010110101010010101011010101001100110011001100110011001100110,
64'b0110100110010110011010011001011010010110100101101001011010010110,
64'b0110100101101001100101101001011001100110100110011001100101100110,
64'b1100110011001100110011001100110001100110100110011001100101100110,
64'b0110011001100110011001100110011011111111000000001111111100000000,
64'b0101101001011010010110100101101000110011110011000011001111001100,
64'b1010101001010101010101011010101001101001011010011001011010010110,
64'b1111111100000000111111110000000001011010010110100101101001011010,
64'b0011001100110011110011001100110011110000111100001111000011110000,
64'b0101010101010101101010101010101011000011001111001100001100111100,
64'b1001011010010110100101101001011011111111000000001111111100000000,
64'b1111111100000000111111110000000001010101010101011010101010101010,
64'b1010101010101010101010101010101000111100001111000011110000111100,
64'b0011001100110011110011001100110000111100001111000011110000111100,
64'b0011110011000011110000110011110011000011001111001100001100111100,
64'b1100001100111100110000110011110011000011110000110011110000111100,
64'b0101101001011010010110100101101001101001011010011001011010010110,
64'b0011110000111100001111000011110001010101010101011010101010101010,
64'b0011001111001100001100111100110000001111000011111111000011110000,
64'b0011001100110011110011001100110011000011001111001100001100111100,
64'b1010101010101010101010101010101010011001011001101001100101100110,
64'b1010101010101010101010101010101011111111000000001111111100000000,
64'b1001100101100110100110010110011011110000000011110000111111110000,
64'b1010101001010101010101011010101011111111111111110000000000000000,
64'b1010101010101010101010101010101011001100110011001100110011001100,
64'b0110100110010110011010011001011010100101010110101010010101011010,
64'b1111000000001111000011111111000000001111111100000000111111110000,
64'b0011001100110011110011001100110011110000000011110000111111110000,
64'b0110100101101001100101101001011000001111111100000000111111110000,
64'b1001011010010110100101101001011001101001100101100110100110010110,
64'b1100110000110011001100111100110001100110011001100110011001100110,
64'b1100001100111100110000110011110001010101101010100101010110101010,
64'b1010101010101010101010101010101001011010101001011010010101011010,
64'b1001100101100110100110010110011000111100001111000011110000111100,
64'b0011110000111100001111000011110011111111111111110000000000000000,
64'b0011110011000011110000110011110000000000111111111111111100000000,
64'b1111000011110000111100001111000010101010101010101010101010101010,
64'b0011001100110011110011001100110001011010010110100101101001011010,
64'b1001100110011001011001100110011011001100001100110011001111001100,
64'b0000000000000000000000000000000000000000111111111111111100000000,
64'b0011001111001100001100111100110000000000111111111111111100000000,
64'b0101101001011010010110100101101010101010010101010101010110101010,
64'b1100110011001100110011001100110000111100110000111100001100111100,
64'b1100110011001100110011001100110000111100001111000011110000111100,
64'b1001011010010110100101101001011000110011001100111100110011001100,
64'b1001011010010110100101101001011011001100001100110011001111001100,
64'b1100001100111100110000110011110010100101010110101010010101011010,
64'b0000111111110000000011111111000011110000111100001111000011110000,
64'b1111000000001111000011111111000010101010010101010101010110101010,
64'b0101010110101010010101011010101010100101101001010101101001011010,
64'b1111000011110000111100001111000001100110100110011001100101100110,
64'b1001011010010110100101101001011010101010010101010101010110101010,
64'b1010101010101010101010101010101001010101101010100101010110101010,
64'b0000111100001111111100001111000000111100110000111100001100111100,
64'b0011001111001100001100111100110010101010010101010101010110101010,
64'b1111000011110000111100001111000011111111111111110000000000000000,
64'b1111000011110000111100001111000001100110100110011001100101100110,
64'b1100001100111100110000110011110000111100110000111100001100111100,
64'b1100001100111100110000110011110011111111111111110000000000000000,
64'b0000111111110000000011111111000001100110011001100110011001100110,
64'b1111000000001111000011111111000000001111111100000000111111110000,
64'b1111111111111111000000000000000011001100001100110011001111001100,
64'b0101101001011010010110100101101001011010101001011010010101011010,
64'b1010101001010101010101011010101000111100001111000011110000111100,
64'b0110011001100110011001100110011000111100110000111100001100111100,
64'b1100110000110011001100111100110010011001011001101001100101100110,
64'b1001011010010110100101101001011010011001100110010110011001100110,
64'b1001011001101001011010011001011010101010010101010101010110101010,
64'b0101101001011010010110100101101000001111111100000000111111110000,
64'b0011110011000011110000110011110010101010101010101010101010101010,
64'b0011110000111100001111000011110010010110100101101001011010010110,
64'b1010101001010101010101011010101011110000111100001111000011110000,
64'b0000000000000000000000000000000001101001100101100110100110010110,
64'b1111000000001111000011111111000000000000111111111111111100000000,
64'b0101010110101010010101011010101000001111000011111111000011110000,
64'b0101101010100101101001010101101001100110100110011001100101100110,
64'b0110011001100110011001100110011010100101010110101010010101011010,
64'b0011001111001100001100111100110011110000000011110000111111110000,
64'b0000111111110000000011111111000001101001011010011001011010010110,
64'b0000000000000000000000000000000000111100001111000011110000111100,
64'b0000111100001111111100001111000010011001100110010110011001100110,
64'b0011110000111100001111000011110010101010010101010101010110101010,
64'b0011001111001100001100111100110011001100110011001100110011001100,
64'b0110100101101001100101101001011011000011001111001100001100111100,
64'b0110100101101001100101101001011011111111000000001111111100000000,
64'b0101010110101010010101011010101011000011001111001100001100111100,
64'b1010101001010101010101011010101011111111111111110000000000000000,
64'b1001100110011001011001100110011001010101101010100101010110101010,
64'b1100110000110011001100111100110001101001011010011001011010010110,
64'b1001011010010110100101101001011001100110100110011001100101100110,
64'b0000111100001111111100001111000000000000111111111111111100000000,
64'b0000000011111111111111110000000001101001100101100110100110010110,
64'b0000000000000000000000000000000010100101010110101010010101011010,
64'b1111111100000000111111110000000000111100001111000011110000111100,
64'b1010010101011010101001010101101010011001100110010110011001100110,
64'b0000111100001111111100001111000001011010010110100101101001011010,
64'b1100001100111100110000110011110011110000000011110000111111110000,
64'b0110100110010110011010011001011011111111111111110000000000000000,
64'b0110011001100110011001100110011000001111111100000000111111110000,
64'b0110100101101001100101101001011011110000111100001111000011110000,
64'b0110100110010110011010011001011001100110100110011001100101100110,
64'b0110011001100110011001100110011000000000111111111111111100000000,
64'b0011110011000011110000110011110000111100001111000011110000111100,
64'b0101101001011010010110100101101011110000000011110000111111110000,
64'b0101010110101010010101011010101010010110100101101001011010010110,
64'b1100001100111100110000110011110010100101101001010101101001011010,
64'b1100110000110011001100111100110000111100001111000011110000111100,
64'b0110100101101001100101101001011010011001011001101001100101100110,
64'b0011110011000011110000110011110001011010101001011010010101011010,
64'b1001011010010110100101101001011011001100110011001100110011001100,
64'b0110011010011001100110010110011011110000111100001111000011110000,
64'b1100001100111100110000110011110010101010101010101010101010101010,
64'b1001100101100110100110010110011011111111000000001111111100000000,
64'b0110100101101001100101101001011011000011110000110011110000111100,
64'b1111111111111111000000000000000001010101010101011010101010101010,
64'b1010010101011010101001010101101010100101010110101010010101011010,
64'b0011110000111100001111000011110000000000111111111111111100000000,
64'b0011001111001100001100111100110001101001100101100110100110010110,
64'b1001100110011001011001100110011000110011110011000011001111001100,
64'b0011110011000011110000110011110010100101010110101010010101011010,
64'b1100110011001100110011001100110011000011110000110011110000111100,
64'b1001100101100110100110010110011011001100001100110011001111001100,
64'b1010010110100101010110100101101001011010010110100101101001011010,
64'b1001100110011001011001100110011011111111000000001111111100000000,
64'b0101101001011010010110100101101011001100110011001100110011001100,
64'b1001100110011001011001100110011011111111111111110000000000000000,
64'b0011110000111100001111000011110000001111111100000000111111110000,
64'b0110100101101001100101101001011001100110011001100110011001100110,
64'b0011001111001100001100111100110001100110100110011001100101100110,
64'b1010101010101010101010101010101011111111111111110000000000000000,
64'b0000111111110000000011111111000010010110011010010110100110010110,
64'b0101010110101010010101011010101000001111000011111111000011110000,
64'b0110100101101001100101101001011011001100001100110011001111001100,
64'b1111111100000000111111110000000000001111111100000000111111110000,
64'b0000000000000000000000000000000010100101101001010101101001011010,
64'b1111111111111111000000000000000010011001011001101001100101100110,
64'b1100110011001100110011001100110011111111111111110000000000000000,
64'b0110011001100110011001100110011011110000111100001111000011110000,
64'b1001011010010110100101101001011000000000000000000000000000000000,
64'b1010010101011010101001010101101010101010010101010101010110101010,
64'b1100001100111100110000110011110000111100001111000011110000111100,
64'b1010010110100101010110100101101011000011110000110011110000111100,
64'b1100110011001100110011001100110010101010101010101010101010101010,
64'b0000000011111111111111110000000010010110011010010110100110010110,
64'b0011001100110011110011001100110001010101101010100101010110101010,
64'b1100001100111100110000110011110010100101101001010101101001011010,
64'b0101010101010101101010101010101010101010010101010101010110101010,
64'b0000000000000000000000000000000000110011110011000011001111001100,
64'b0000000000000000000000000000000001101001011010011001011010010110,
64'b0101101001011010010110100101101000000000000000000000000000000000,
64'b0011110000111100001111000011110001010101101010100101010110101010,
64'b0110100110010110011010011001011010101010101010101010101010101010,
64'b1100110000110011001100111100110000110011001100111100110011001100,
64'b1111000000001111000011111111000010100101010110101010010101011010,
64'b0011001111001100001100111100110000001111111100000000111111110000,
64'b0101101001011010010110100101101001100110011001100110011001100110,
64'b1111111111111111000000000000000000111100110000111100001100111100,
64'b0101101001011010010110100101101010011001100110010110011001100110,
64'b0101101010100101101001010101101000110011110011000011001111001100,
64'b1100110011001100110011001100110010011001100110010110011001100110,
64'b1010101010101010101010101010101010100101101001010101101001011010,
64'b0000000000000000000000000000000011000011001111001100001100111100,
64'b0011001111001100001100111100110010101010101010101010101010101010,
64'b0000111111110000000011111111000011001100110011001100110011001100,
64'b0011110011000011110000110011110011001100110011001100110011001100,
64'b0000111100001111111100001111000011110000111100001111000011110000,
64'b1010101001010101010101011010101001100110100110011001100101100110,
64'b1010010110100101010110100101101000000000111111111111111100000000,
64'b0011001111001100001100111100110000111100001111000011110000111100,
64'b0000000000000000000000000000000011110000000011110000111111110000,
64'b1001100101100110100110010110011010010110100101101001011010010110,
64'b1100110000110011001100111100110010100101101001010101101001011010,
64'b0101101001011010010110100101101000111100001111000011110000111100,
64'b1100110011001100110011001100110010011001011001101001100101100110,
64'b0000000000000000000000000000000001011010101001011010010101011010,
64'b0000111100001111111100001111000011001100110011001100110011001100,
64'b1111111100000000111111110000000011110000111100001111000011110000,
64'b1111000011110000111100001111000010010110100101101001011010010110,
64'b0011110000111100001111000011110001011010101001011010010101011010,
64'b0110100110010110011010011001011000111100001111000011110000111100,
64'b1111000011110000111100001111000001100110011001100110011001100110,
64'b1100110000110011001100111100110010011001011001101001100101100110,
64'b1001011001101001011010011001011011111111111111110000000000000000,
64'b0011110011000011110000110011110000000000000000000000000000000000,
64'b0110011010011001100110010110011000001111111100000000111111110000,
64'b1100001111000011001111000011110000111100110000111100001100111100,
64'b1100110000110011001100111100110010100101101001010101101001011010,
64'b1111111111111111000000000000000001100110100110011001100101100110,
64'b0011001111001100001100111100110001101001011010011001011010010110,
64'b0011110000111100001111000011110000000000000000000000000000000000,
64'b1010010101011010101001010101101001101001100101100110100110010110,
64'b0011001111001100001100111100110011001100001100110011001111001100,
64'b0101010101010101101010101010101010100101010110101010010101011010,
64'b0000111111110000000011111111000000111100001111000011110000111100,
64'b1100001100111100110000110011110011000011110000110011110000111100,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0110011001100110011001100110011010101010101010101010101010101010,
64'b0000111111110000000011111111000000000000111111111111111100000000,
64'b0110011010011001100110010110011011110000000011110000111111110000,
64'b0110100110010110011010011001011010011001011001101001100101100110,
64'b0101010101010101101010101010101001101001011010011001011010010110,
64'b1001011001101001011010011001011001101001100101100110100110010110,
64'b0011001111001100001100111100110010101010101010101010101010101010,
64'b1001011001101001011010011001011000111100110000111100001100111100,
64'b0011001100110011110011001100110000001111000011111111000011110000,
64'b1010010101011010101001010101101001100110100110011001100101100110,
64'b0101101010100101101001010101101000001111111100000000111111110000,
64'b0011110000111100001111000011110000001111111100000000111111110000,
64'b1001011001101001011010011001011010101010101010101010101010101010,
64'b0000000011111111111111110000000011001100110011001100110011001100,
64'b0110011001100110011001100110011011111111111111110000000000000000,
64'b0000000000000000000000000000000010101010010101010101010110101010,
64'b0101101001011010010110100101101001101001011010011001011010010110,
64'b0011001100110011110011001100110011000011001111001100001100111100,
64'b1010010110100101010110100101101010010110011010010110100110010110,
64'b0110011001100110011001100110011011001100110011001100110011001100,
64'b1001011001101001011010011001011011110000000011110000111111110000,
64'b0101101001011010010110100101101001010101101010100101010110101010,
64'b0110011010011001100110010110011001101001011010011001011010010110,
64'b1100110000110011001100111100110010101010010101010101010110101010,
64'b1010010101011010101001010101101000000000111111111111111100000000,
64'b0011110011000011110000110011110011001100110011001100110011001100,
64'b0101010101010101101010101010101011110000111100001111000011110000,
64'b1001011010010110100101101001011000000000000000000000000000000000,
64'b0000000000000000000000000000000010011001100110010110011001100110,
64'b0011001111001100001100111100110001101001100101100110100110010110,
64'b1111000011110000111100001111000001011010101001011010010101011010,
64'b1001100101100110100110010110011000111100110000111100001100111100,
64'b1001011010010110100101101001011001011010010110100101101001011010,
64'b1100110000110011001100111100110010101010010101010101010110101010,
64'b1010010101011010101001010101101010011001100110010110011001100110,
64'b1010101001010101010101011010101011000011001111001100001100111100,
64'b0101010101010101101010101010101010011001100110010110011001100110,
64'b1010101010101010101010101010101001010101010101011010101010101010,
64'b0110011001100110011001100110011001011010010110100101101001011010,
64'b0101101010100101101001010101101011111111000000001111111100000000,
64'b0000111100001111111100001111000000000000000000000000000000000000,
64'b1100001111000011001111000011110000111100001111000011110000111100,
64'b1100001100111100110000110011110010010110011010010110100110010110,
64'b0000000011111111111111110000000011001100001100110011001111001100,
64'b1111000000001111000011111111000001011010101001011010010101011010,
64'b1111111100000000111111110000000010011001011001101001100101100110,
64'b0101010101010101101010101010101000110011001100111100110011001100,
64'b0101101010100101101001010101101010010110100101101001011010010110,
64'b0101101010100101101001010101101001011010101001011010010101011010,
64'b1001011010010110100101101001011000111100001111000011110000111100,
64'b1010101001010101010101011010101001100110011001100110011001100110,
64'b1010101001010101010101011010101010011001011001101001100101100110,
64'b1111000011110000111100001111000011111111111111110000000000000000,
64'b0011001100110011110011001100110000000000000000000000000000000000,
64'b0110011010011001100110010110011000001111111100000000111111110000,
64'b1001011010010110100101101001011000111100110000111100001100111100,
64'b0000000000000000000000000000000010100101101001010101101001011010,
64'b1001100110011001011001100110011001100110100110011001100101100110,
64'b1001011010010110100101101001011010010110100101101001011010010110,
64'b0110011001100110011001100110011010101010101010101010101010101010,
64'b0110011010011001100110010110011001010101101010100101010110101010,
64'b0110011010011001100110010110011010100101101001010101101001011010,
64'b0110100110010110011010011001011001010101101010100101010110101010,
64'b0011001100110011110011001100110011110000000011110000111111110000,
64'b1001100110011001011001100110011001010101101010100101010110101010,
64'b0101010110101010010101011010101000111100110000111100001100111100,
64'b1111000011110000111100001111000011001100001100110011001111001100,
64'b0110100101101001100101101001011011000011001111001100001100111100,
64'b0110100110010110011010011001011000111100001111000011110000111100,
64'b0000000000000000000000000000000001100110100110011001100101100110,
64'b0011110000111100001111000011110001011010101001011010010101011010,
64'b0110100110010110011010011001011001010101101010100101010110101010,
64'b0110011001100110011001100110011000111100001111000011110000111100,
64'b1111111111111111000000000000000000001111000011111111000011110000,
64'b0000000011111111111111110000000001011010010110100101101001011010,
64'b0110011010011001100110010110011001101001011010011001011010010110,
64'b0011110011000011110000110011110011001100110011001100110011001100,
64'b0000000011111111111111110000000000001111111100000000111111110000,
64'b1010010101011010101001010101101011001100110011001100110011001100,
64'b1001100110011001011001100110011011000011001111001100001100111100,
64'b0000000011111111111111110000000010011001011001101001100101100110,
64'b0101101001011010010110100101101011000011110000110011110000111100,
64'b1111111111111111000000000000000000111100001111000011110000111100,
64'b0011110000111100001111000011110001010101010101011010101010101010,
64'b1111111100000000111111110000000001011010010110100101101001011010,
64'b1100110011001100110011001100110010100101010110101010010101011010,
64'b0011110000111100001111000011110011111111000000001111111100000000,
64'b0011110011000011110000110011110010011001011001101001100101100110,
64'b1001100110011001011001100110011011000011001111001100001100111100,
64'b1001011010010110100101101001011001011010010110100101101001011010,
64'b1100001100111100110000110011110000000000111111111111111100000000,
64'b0101101001011010010110100101101011110000111100001111000011110000,
64'b0101101010100101101001010101101011110000000011110000111111110000,
64'b1001011010010110100101101001011011000011110000110011110000111100,
64'b0101010101010101101010101010101000001111111100000000111111110000,
64'b1111111111111111000000000000000010100101010110101010010101011010,
64'b1001011010010110100101101001011011001100110011001100110011001100,
64'b0011110000111100001111000011110010011001011001101001100101100110,
64'b0101101001011010010110100101101001100110100110011001100101100110,
64'b0000111111110000000011111111000011111111111111110000000000000000,
64'b1111000000001111000011111111000011000011110000110011110000111100,
64'b1001011010010110100101101001011011110000000011110000111111110000,
64'b0110100110010110011010011001011000110011110011000011001111001100,
64'b1111000000001111000011111111000011111111111111110000000000000000,
64'b0011001111001100001100111100110001010101101010100101010110101010,
64'b1100110000110011001100111100110000000000111111111111111100000000,
64'b0110100110010110011010011001011010100101010110101010010101011010,
64'b1100110011001100110011001100110010101010010101010101010110101010,
64'b1010101010101010101010101010101011001100001100110011001111001100,
64'b0110100110010110011010011001011011110000111100001111000011110000,
64'b0000111111110000000011111111000000111100001111000011110000111100,
64'b1100001100111100110000110011110010011001100110010110011001100110,
64'b0011110011000011110000110011110010010110100101101001011010010110,
64'b0110100101101001100101101001011011001100110011001100110011001100,
64'b1001100101100110100110010110011001011010101001011010010101011010,
64'b1111000011110000111100001111000001101001100101100110100110010110,
64'b1001011010010110100101101001011010010110011010010110100110010110,
64'b1001100101100110100110010110011010100101010110101010010101011010,
64'b0110100110010110011010011001011010011001011001101001100101100110,
64'b0101010110101010010101011010101010100101010110101010010101011010,
64'b0011110011000011110000110011110011111111000000001111111100000000,
64'b0011001100110011110011001100110001011010010110100101101001011010,
64'b0000111100001111111100001111000001100110011001100110011001100110,
64'b1100001100111100110000110011110000110011110011000011001111001100,
64'b1010101001010101010101011010101000111100001111000011110000111100,
64'b1100110000110011001100111100110001101001100101100110100110010110,
64'b0000000000000000000000000000000011110000111100001111000011110000,
64'b1001100110011001011001100110011011001100001100110011001111001100,
64'b0011001100110011110011001100110010010110011010010110100110010110,
64'b0101010101010101101010101010101000111100110000111100001100111100,
64'b1111111100000000111111110000000001100110100110011001100101100110,
64'b0101101001011010010110100101101011000011110000110011110000111100,
64'b1111000011110000111100001111000011001100001100110011001111001100,
64'b0011110000111100001111000011110011111111111111110000000000000000,
64'b1010010110100101010110100101101000110011110011000011001111001100,
64'b0110011001100110011001100110011000111100001111000011110000111100,
64'b1001100101100110100110010110011011110000111100001111000011110000,
64'b1100001111000011001111000011110000001111111100000000111111110000,
64'b1001100110011001011001100110011000111100110000111100001100111100,
64'b1100001100111100110000110011110011111111000000001111111100000000,
64'b1100110011001100110011001100110000001111000011111111000011110000,
64'b1001011001101001011010011001011010010110011010010110100110010110,
64'b1111000000001111000011111111000001011010101001011010010101011010,
64'b0110100110010110011010011001011001101001011010011001011010010110,
64'b0101010101010101101010101010101010100101010110101010010101011010,
64'b0011110011000011110000110011110010100101101001010101101001011010,
64'b1100001111000011001111000011110010101010101010101010101010101010,
64'b1100110000110011001100111100110010100101101001010101101001011010,
64'b1010010101011010101001010101101000001111111100000000111111110000,
64'b0000000000000000000000000000000011111111000000001111111100000000,
64'b0000111111110000000011111111000000000000111111111111111100000000,
64'b1001011010010110100101101001011011110000000011110000111111110000,
64'b0101101010100101101001010101101001010101010101011010101010101010,
64'b1111000011110000111100001111000011111111000000001111111100000000,
64'b0011110011000011110000110011110010010110011010010110100110010110,
64'b1010101001010101010101011010101001100110100110011001100101100110,
64'b1001011001101001011010011001011001101001100101100110100110010110,
64'b1100110011001100110011001100110001100110100110011001100101100110,
64'b0101101010100101101001010101101000110011110011000011001111001100,
64'b1010010101011010101001010101101001100110011001100110011001100110,
64'b1010010110100101010110100101101000110011110011000011001111001100,
64'b0110011010011001100110010110011010101010010101010101010110101010,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000011111111111111110000000001010101010101011010101010101010,
64'b1100001100111100110000110011110010101010010101010101010110101010,
64'b1100110000110011001100111100110001100110011001100110011001100110,
64'b0101010110101010010101011010101001010101010101011010101010101010,
64'b1111000000001111000011111111000000111100110000111100001100111100,
64'b1001100110011001011001100110011001101001011010011001011010010110,
64'b1001011001101001011010011001011010010110011010010110100110010110,
64'b0101101001011010010110100101101011000011110000110011110000111100,
64'b1100110000110011001100111100110010100101101001010101101001011010,
64'b0110011010011001100110010110011000111100001111000011110000111100,
64'b0011001111001100001100111100110000001111000011111111000011110000,
64'b0110100101101001100101101001011000110011001100111100110011001100,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b0101010101010101101010101010101011001100110011001100110011001100,
64'b0101101010100101101001010101101010011001100110010110011001100110,
64'b0000111100001111111100001111000010010110100101101001011010010110,
64'b1001100110011001011001100110011011001100110011001100110011001100,
64'b0000000011111111111111110000000001011010101001011010010101011010,
64'b1001011010010110100101101001011001101001100101100110100110010110,
64'b1001011001101001011010011001011010010110011010010110100110010110,
64'b1001100101100110100110010110011010100101010110101010010101011010,
64'b0000111100001111111100001111000010011001011001101001100101100110,
64'b0110100101101001100101101001011010100101010110101010010101011010,
64'b1010010110100101010110100101101011111111000000001111111100000000,
64'b1100001100111100110000110011110001011010010110100101101001011010,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b1111111100000000111111110000000000000000111111111111111100000000,
64'b0101101001011010010110100101101000110011001100111100110011001100,
64'b0000111100001111111100001111000001011010010110100101101001011010,
64'b1001011001101001011010011001011001010101101010100101010110101010,
64'b0000111100001111111100001111000001010101101010100101010110101010,
64'b0011001100110011110011001100110000110011110011000011001111001100,
64'b0101010110101010010101011010101010100101010110101010010101011010,
64'b0011001111001100001100111100110010101010010101010101010110101010,
64'b1010010101011010101001010101101010011001011001101001100101100110,
64'b1001011001101001011010011001011011001100110011001100110011001100,
64'b0110100101101001100101101001011000000000000000000000000000000000,
64'b0000000011111111111111110000000001010101101010100101010110101010,
64'b0101010110101010010101011010101000001111111100000000111111110000,
64'b0000000011111111111111110000000011111111111111110000000000000000,
64'b0110100110010110011010011001011001011010010110100101101001011010,
64'b1111000000001111000011111111000010011001011001101001100101100110,
64'b0000000000000000000000000000000000110011001100111100110011001100,
64'b0101101010100101101001010101101000110011001100111100110011001100,
64'b0110100101101001100101101001011000001111000011111111000011110000,
64'b1100110000110011001100111100110011001100001100110011001111001100,
64'b0011110011000011110000110011110000110011001100111100110011001100,
64'b0110100101101001100101101001011001101001011010011001011010010110,
64'b1010101010101010101010101010101011110000111100001111000011110000,
64'b0000000011111111111111110000000000000000000000000000000000000000,
64'b0101010110101010010101011010101000110011001100111100110011001100,
64'b0011001111001100001100111100110011111111000000001111111100000000,
64'b1010101001010101010101011010101000000000000000000000000000000000,
64'b1100110000110011001100111100110010011001011001101001100101100110,
64'b0000111111110000000011111111000011000011110000110011110000111100,
64'b0011110011000011110000110011110011110000111100001111000011110000,
64'b1100001100111100110000110011110001011010010110100101101001011010,
64'b0101101010100101101001010101101001010101101010100101010110101010,
64'b1111000000001111000011111111000010100101101001010101101001011010,
64'b0110100101101001100101101001011001011010010110100101101001011010,
64'b1100110011001100110011001100110001101001100101100110100110010110,
64'b1111000000001111000011111111000001010101101010100101010110101010,
64'b1001011010010110100101101001011000000000000000000000000000000000,
64'b1001100101100110100110010110011011110000111100001111000011110000,
64'b1010010101011010101001010101101010101010101010101010101010101010,
64'b0011001100110011110011001100110000000000000000000000000000000000,
64'b1010010110100101010110100101101011000011110000110011110000111100,
64'b1010101001010101010101011010101000001111111100000000111111110000,
64'b1111000000001111000011111111000001010101101010100101010110101010,
64'b0101101010100101101001010101101000110011110011000011001111001100,
64'b1100110000110011001100111100110000110011001100111100110011001100,
64'b1010101001010101010101011010101000110011110011000011001111001100,
64'b0110100110010110011010011001011010011001011001101001100101100110,
64'b0101101001011010010110100101101000111100110000111100001100111100,
64'b0000000011111111111111110000000000110011001100111100110011001100,
64'b0110100110010110011010011001011000000000000000000000000000000000,
64'b1100001111000011001111000011110011111111000000001111111100000000,
64'b0011001111001100001100111100110011001100110011001100110011001100,
64'b0000111111110000000011111111000000000000000000000000000000000000,
64'b1100001100111100110000110011110000001111111100000000111111110000,
64'b1001011010010110100101101001011010101010010101010101010110101010,
64'b0011110000111100001111000011110000110011001100111100110011001100,
64'b0110100110010110011010011001011000001111000011111111000011110000,
64'b1001011010010110100101101001011011110000111100001111000011110000,
64'b1100110000110011001100111100110010100101101001010101101001011010,
64'b1010010110100101010110100101101011000011110000110011110000111100,
64'b1001011010010110100101101001011011110000000011110000111111110000,
64'b0110100110010110011010011001011001011010010110100101101001011010,
64'b1111111100000000111111110000000010101010101010101010101010101010,
64'b0000111100001111111100001111000011111111111111110000000000000000,
64'b0000111111110000000011111111000011110000111100001111000011110000,
64'b0101010101010101101010101010101010101010101010101010101010101010,
64'b1010101001010101010101011010101000000000111111111111111100000000,
64'b1100110000110011001100111100110000110011001100111100110011001100,
64'b1001100110011001011001100110011001011010010110100101101001011010,
64'b0011001111001100001100111100110001010101101010100101010110101010,
64'b1111000000001111000011111111000001010101101010100101010110101010,
64'b0101101010100101101001010101101000110011110011000011001111001100,
64'b1010101010101010101010101010101010100101010110101010010101011010,
64'b1100110011001100110011001100110010101010010101010101010110101010,
64'b1010101010101010101010101010101010011001011001101001100101100110,
64'b1001011010010110100101101001011011001100110011001100110011001100,
64'b1111111111111111000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000001010101101010100101010110101010,
64'b1100110011001100110011001100110000110011110011000011001111001100,
64'b1001100110011001011001100110011010100101101001010101101001011010,
64'b1010010110100101010110100101101001010101010101011010101010101010,
64'b1001011010010110100101101001011000001111000011111111000011110000,
64'b1010010110100101010110100101101000111100001111000011110000111100,
64'b0000000011111111111111110000000000000000000000000000000000000000,
64'b0110011010011001100110010110011001011010101001011010010101011010,
64'b0110011001100110011001100110011011111111111111110000000000000000,
64'b1111000011110000111100001111000010010110011010010110100110010110,
64'b1100110011001100110011001100110011111111000000001111111100000000,
64'b1100001100111100110000110011110010011001100110010110011001100110,
64'b0000000000000000000000000000000000000000111111111111111100000000,
64'b1010101010101010101010101010101010011001011001101001100101100110,
64'b1010010101011010101001010101101001011010101001011010010101011010,
64'b0110011001100110011001100110011001101001100101100110100110010110,
64'b1001011001101001011010011001011001101001011010011001011010010110,
64'b1111111111111111000000000000000011000011110000110011110000111100,
64'b0011110011000011110000110011110010101010010101010101010110101010,
64'b0110011001100110011001100110011000110011001100111100110011001100,
64'b0011110011000011110000110011110010011001100110010110011001100110,
64'b1010010101011010101001010101101010011001011001101001100101100110,
64'b0101101001011010010110100101101000110011001100111100110011001100,
64'b0110011010011001100110010110011011000011001111001100001100111100,
64'b1001100101100110100110010110011001010101010101011010101010101010,
64'b0000000011111111111111110000000001010101101010100101010110101010,
64'b1001100101100110100110010110011011000011001111001100001100111100,
64'b1001100110011001011001100110011011001100001100110011001111001100,
64'b0110011001100110011001100110011010010110011010010110100110010110,
64'b0011001111001100001100111100110011000011001111001100001100111100,
64'b0011110011000011110000110011110010100101010110101010010101011010,
64'b0101010110101010010101011010101010011001100110010110011001100110,
64'b1010010110100101010110100101101001011010010110100101101001011010,
64'b1010010110100101010110100101101010010110100101101001011010010110,
64'b0101010101010101101010101010101001101001011010011001011010010110,
64'b1001011010010110100101101001011011110000111100001111000011110000,
64'b0101010110101010010101011010101001011010101001011010010101011010,
64'b0000000000000000000000000000000011001100110011001100110011001100,
64'b1111111100000000111111110000000010011001100110010110011001100110,
64'b1100001100111100110000110011110000001111111100000000111111110000,
64'b0011110000111100001111000011110010100101101001010101101001011010,
64'b1001011010010110100101101001011010010110011010010110100110010110,
64'b0000111100001111111100001111000001011010101001011010010101011010,
64'b1111000000001111000011111111000011001100001100110011001111001100,
64'b1001100110011001011001100110011000111100001111000011110000111100,
64'b0011001111001100001100111100110010011001011001101001100101100110,
64'b1001100101100110100110010110011011000011001111001100001100111100,
64'b0110011001100110011001100110011011000011001111001100001100111100,
64'b0110100110010110011010011001011001010101101010100101010110101010,
64'b0011001100110011110011001100110011001100001100110011001111001100,
64'b0000000000000000000000000000000001011010010110100101101001011010,
64'b1111111111111111000000000000000000111100001111000011110000111100,
64'b0000111111110000000011111111000001010101101010100101010110101010,
64'b0101101001011010010110100101101011001100110011001100110011001100,
64'b1001100101100110100110010110011011001100001100110011001111001100,
64'b1111000000001111000011111111000001101001100101100110100110010110,
64'b0011110000111100001111000011110000110011110011000011001111001100,
64'b1001100110011001011001100110011010101010010101010101010110101010,
64'b1001011010010110100101101001011011110000111100001111000011110000,
64'b1001011001101001011010011001011010100101101001010101101001011010,
64'b0000111111110000000011111111000011000011110000110011110000111100,
64'b1001100110011001011001100110011010010110011010010110100110010110,
64'b0110011010011001100110010110011010011001011001101001100101100110,
64'b1100001111000011001111000011110011110000000011110000111111110000,
64'b0000000011111111111111110000000000001111000011111111000011110000,
64'b0000000000000000000000000000000010011001011001101001100101100110,
64'b0110011001100110011001100110011001011010010110100101101001011010,
64'b1001100110011001011001100110011000001111000011111111000011110000,
64'b0000111111110000000011111111000010010110011010010110100110010110,
64'b0011001100110011110011001100110000001111000011111111000011110000,
64'b0011001100110011110011001100110000110011001100111100110011001100,
64'b0101101010100101101001010101101001010101101010100101010110101010,
64'b0110100101101001100101101001011000110011110011000011001111001100,
64'b1001100110011001011001100110011010100101010110101010010101011010,
64'b1001100101100110100110010110011010010110011010010110100110010110,
64'b1111111100000000111111110000000001101001011010011001011010010110,
64'b1100110000110011001100111100110000000000111111111111111100000000,
64'b0101010110101010010101011010101001010101101010100101010110101010,
64'b1111111100000000111111110000000010010110100101101001011010010110,
64'b0110100110010110011010011001011000110011110011000011001111001100,
64'b0110011001100110011001100110011011111111000000001111111100000000,
64'b1010010101011010101001010101101010010110011010010110100110010110,
64'b0110011010011001100110010110011001010101101010100101010110101010,
64'b0101010101010101101010101010101001011010010110100101101001011010,
64'b0101010110101010010101011010101010011001100110010110011001100110,
64'b0011110000111100001111000011110000001111000011111111000011110000,
64'b1010010101011010101001010101101011001100001100110011001111001100,
64'b1100110000110011001100111100110000111100110000111100001100111100,
64'b0110100110010110011010011001011001101001100101100110100110010110,
64'b0110011001100110011001100110011001010101010101011010101010101010,
64'b1001100101100110100110010110011010011001100110010110011001100110,
64'b0101010110101010010101011010101011000011001111001100001100111100,
64'b0011110011000011110000110011110010100101101001010101101001011010,
64'b0011110000111100001111000011110011111111111111110000000000000000,
64'b1100110000110011001100111100110000111100110000111100001100111100,
64'b1100001111000011001111000011110010011001100110010110011001100110,
64'b0110011001100110011001100110011000110011110011000011001111001100,
64'b1001100110011001011001100110011000111100001111000011110000111100,
64'b0000111111110000000011111111000001010101101010100101010110101010,
64'b1100110000110011001100111100110010100101101001010101101001011010,
64'b0000111100001111111100001111000001011010101001011010010101011010,
64'b1001011001101001011010011001011010010110011010010110100110010110,
64'b0011110000111100001111000011110011001100110011001100110011001100,
64'b1100001111000011001111000011110010010110100101101001011010010110,
64'b1100110011001100110011001100110010100101010110101010010101011010,
64'b1111000000001111000011111111000000110011110011000011001111001100,
64'b1010010101011010101001010101101010101010101010101010101010101010,
64'b0000111100001111111100001111000001011010101001011010010101011010,
64'b1010010101011010101001010101101010010110100101101001011010010110,
64'b1001011010010110100101101001011010100101101001010101101001011010,
64'b0011110000111100001111000011110000001111111100000000111111110000,
64'b1010101001010101010101011010101000110011001100111100110011001100,
64'b0000111100001111111100001111000000110011110011000011001111001100,
64'b0101010110101010010101011010101001100110100110011001100101100110,
64'b1001011001101001011010011001011010010110011010010110100110010110,
64'b1010010101011010101001010101101001011010010110100101101001011010,
64'b0000111111110000000011111111000011000011001111001100001100111100,
64'b0101101001011010010110100101101000110011110011000011001111001100,
64'b0000000011111111111111110000000000001111000011111111000011110000,
64'b0110011010011001100110010110011011001100110011001100110011001100,
64'b1111111100000000111111110000000011001100001100110011001111001100,
64'b0110011010011001100110010110011001101001100101100110100110010110,
64'b1100001100111100110000110011110000110011110011000011001111001100,
64'b0000111111110000000011111111000010101010010101010101010110101010,
64'b0011001100110011110011001100110011110000111100001111000011110000,
64'b0101010110101010010101011010101010100101101001010101101001011010,
64'b1001100110011001011001100110011011000011110000110011110000111100,
64'b0011110011000011110000110011110010010110011010010110100110010110,
64'b0110011010011001100110010110011010011001011001101001100101100110,
64'b0000000011111111111111110000000011110000000011110000111111110000,
64'b0011001111001100001100111100110011110000111100001111000011110000,
64'b1100001100111100110000110011110001101001011010011001011010010110,
64'b0110011001100110011001100110011000000000111111111111111100000000,
64'b1100001100111100110000110011110011110000000011110000111111110000,
64'b0101010101010101101010101010101000110011110011000011001111001100,
64'b0011001111001100001100111100110010100101010110101010010101011010,
64'b1010010110100101010110100101101010101010101010101010101010101010,
64'b0000000000000000000000000000000011000011001111001100001100111100,
64'b1111000011110000111100001111000010010110011010010110100110010110,
64'b0011001111001100001100111100110000110011001100111100110011001100,
64'b1100001100111100110000110011110010010110011010010110100110010110,
64'b1010010101011010101001010101101010100101010110101010010101011010,
64'b0011110000111100001111000011110010100101101001010101101001011010,
64'b1111111100000000111111110000000011000011001111001100001100111100,
64'b1001100110011001011001100110011001101001100101100110100110010110,
64'b0101101001011010010110100101101001010101010101011010101010101010,
64'b0011001100110011110011001100110010101010010101010101010110101010,
64'b1001100110011001011001100110011010100101101001010101101001011010,
64'b1001011001101001011010011001011011001100001100110011001111001100,
64'b1001011001101001011010011001011011001100110011001100110011001100,
64'b1010101010101010101010101010101011110000000011110000111111110000,
64'b0000111111110000000011111111000000111100110000111100001100111100,
64'b0011110011000011110000110011110001011010010110100101101001011010,
64'b0011001100110011110011001100110010010110011010010110100110010110,
64'b0110100101101001100101101001011001100110100110011001100101100110,
64'b0011001111001100001100111100110000110011110011000011001111001100,
64'b1111111100000000111111110000000010100101010110101010010101011010,
64'b0101010110101010010101011010101010010110011010010110100110010110,
64'b1111111100000000111111110000000011001100110011001100110011001100,
64'b0011001111001100001100111100110010011001100110010110011001100110,
64'b1100001111000011001111000011110010011001011001101001100101100110,
64'b1010010110100101010110100101101010100101101001010101101001011010,
64'b0011001111001100001100111100110001011010010110100101101001011010,
64'b0110011001100110011001100110011000000000111111111111111100000000,
64'b1111000000001111000011111111000001011010101001011010010101011010,
64'b1100001111000011001111000011110010011001011001101001100101100110,
64'b1001100101100110100110010110011000111100110000111100001100111100,
64'b1100110011001100110011001100110001101001011010011001011010010110,
64'b1001100110011001011001100110011010100101101001010101101001011010,
64'b1111111100000000111111110000000000110011110011000011001111001100,
64'b1001100110011001011001100110011000111100110000111100001100111100,
64'b1111111111111111000000000000000001011010010110100101101001011010,
64'b0000111100001111111100001111000000111100001111000011110000111100,
64'b0000111111110000000011111111000001101001011010011001011010010110,
64'b1001100101100110100110010110011000110011110011000011001111001100,
64'b1010010110100101010110100101101010011001011001101001100101100110,
64'b0011110000111100001111000011110011111111111111110000000000000000,
64'b0000000011111111111111110000000001100110100110011001100101100110,
64'b1010010101011010101001010101101001101001011010011001011010010110,
64'b0110100101101001100101101001011011110000000011110000111111110000,
64'b1111000011110000111100001111000001101001100101100110100110010110,
64'b0011110000111100001111000011110010011001011001101001100101100110,
64'b1010101010101010101010101010101001011010010110100101101001011010,
64'b0101010110101010010101011010101011110000000011110000111111110000,
64'b1100110011001100110011001100110010011001011001101001100101100110,
64'b1001011010010110100101101001011000001111111100000000111111110000,
64'b1111111100000000111111110000000011000011001111001100001100111100,
64'b1111000000001111000011111111000010100101101001010101101001011010,
64'b1001011001101001011010011001011011000011110000110011110000111100,
64'b1010010101011010101001010101101000000000000000000000000000000000,
64'b0000111100001111111100001111000001101001011010011001011010010110,
64'b0101010101010101101010101010101001101001100101100110100110010110,
64'b0000000000000000000000000000000010101010010101010101010110101010,
64'b1111000011110000111100001111000010010110011010010110100110010110,
64'b0011001111001100001100111100110011000011110000110011110000111100,
64'b0011001111001100001100111100110000110011110011000011001111001100,
64'b0101101010100101101001010101101000000000111111111111111100000000,
64'b1001011010010110100101101001011001101001011010011001011010010110,
64'b0000000000000000000000000000000000000000111111111111111100000000,
64'b1010101010101010101010101010101011110000000011110000111111110000,
64'b0011001100110011110011001100110000110011110011000011001111001100,
64'b0011001111001100001100111100110010100101010110101010010101011010,
64'b0110011010011001100110010110011010101010101010101010101010101010,
64'b0000111111110000000011111111000011000011001111001100001100111100,
64'b0101010110101010010101011010101010010110011010010110100110010110,
64'b0110100110010110011010011001011000110011001100111100110011001100,
64'b0101101001011010010110100101101010010110011010010110100110010110,
64'b0011001100110011110011001100110010100101010110101010010101011010,
64'b0000111111110000000011111111000001011010010110100101101001011010,
64'b1100110000110011001100111100110010010110011010010110100110010110,
64'b0110100110010110011010011001011000001111111100000000111111110000,
64'b0000000000000000000000000000000010010110011010010110100110010110,
64'b1100110011001100110011001100110011111111000000001111111100000000,
64'b1111000011110000111100001111000010010110011010010110100110010110,
64'b1010010110100101010110100101101001101001100101100110100110010110,
64'b1100001111000011001111000011110011001100110011001100110011001100,
64'b1010101001010101010101011010101000000000111111111111111100000000,
64'b0011001100110011110011001100110000001111000011111111000011110000,
64'b0011110011000011110000110011110010011001011001101001100101100110,
64'b0011001111001100001100111100110000110011001100111100110011001100,
64'b1111000011110000111100001111000001011010101001011010010101011010,
64'b0101010110101010010101011010101011001100110011001100110011001100,
64'b1100110000110011001100111100110001010101010101011010101010101010,
64'b1111000000001111000011111111000011001100001100110011001111001100,
64'b1100001100111100110000110011110011111111111111110000000000000000,
64'b1010010110100101010110100101101000000000000000000000000000000000,
64'b1100110011001100110011001100110000001111000011111111000011110000,
64'b1001011001101001011010011001011000110011110011000011001111001100,
64'b1010010101011010101001010101101011110000111100001111000011110000,
64'b0110100101101001100101101001011000001111000011111111000011110000,
64'b0110100110010110011010011001011001100110011001100110011001100110,
64'b1001100110011001011001100110011010101010010101010101010110101010,
64'b0000000011111111111111110000000001010101101010100101010110101010,
64'b1100001100111100110000110011110001011010101001011010010101011010,
64'b0011001111001100001100111100110010100101010110101010010101011010,
64'b0110011010011001100110010110011001100110011001100110011001100110,
64'b1100110000110011001100111100110010100101101001010101101001011010,
64'b1001100110011001011001100110011010101010101010101010101010101010,
64'b0110011010011001100110010110011010101010101010101010101010101010,
64'b0110100110010110011010011001011011111111000000001111111100000000,
64'b1001100101100110100110010110011010100101101001010101101001011010,
64'b0110011010011001100110010110011011111111000000001111111100000000,
64'b0011001111001100001100111100110011111111000000001111111100000000,
64'b1010010110100101010110100101101010010110100101101001011010010110,
64'b1111111100000000111111110000000000110011001100111100110011001100,
64'b1111000000001111000011111111000010011001100110010110011001100110,
64'b0110011010011001100110010110011011001100001100110011001111001100,
64'b0000111111110000000011111111000010011001011001101001100101100110,
64'b0110100101101001100101101001011010010110100101101001011010010110,
64'b1010010110100101010110100101101000110011110011000011001111001100,
64'b1001011010010110100101101001011001100110011001100110011001100110,
64'b0110100101101001100101101001011011001100110011001100110011001100,
64'b1001011001101001011010011001011011111111111111110000000000000000,
64'b1100001111000011001111000011110000110011110011000011001111001100,
64'b1100001111000011001111000011110001010101010101011010101010101010,
64'b1010010110100101010110100101101011111111111111110000000000000000,
64'b0011001111001100001100111100110011000011001111001100001100111100,
64'b0101010101010101101010101010101011110000111100001111000011110000,
64'b0000000011111111111111110000000010010110100101101001011010010110,
64'b0110100101101001100101101001011010100101101001010101101001011010,
64'b0101010110101010010101011010101010010110100101101001011010010110,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b1111111100000000111111110000000001101001011010011001011010010110,
64'b1010101010101010101010101010101011111111000000001111111100000000,
64'b1001011001101001011010011001011010100101101001010101101001011010,
64'b1010010110100101010110100101101000110011110011000011001111001100,
64'b0000000011111111111111110000000000000000000000000000000000000000,
64'b1010010101011010101001010101101011001100110011001100110011001100,
64'b0110100110010110011010011001011001011010010110100101101001011010,
64'b1001011001101001011010011001011001101001011010011001011010010110,
64'b0000111111110000000011111111000000111100001111000011110000111100,
64'b1111000000001111000011111111000001100110011001100110011001100110,
64'b0101010110101010010101011010101000001111111100000000111111110000,
64'b1001100101100110100110010110011010010110100101101001011010010110,
64'b0000111111110000000011111111000001100110011001100110011001100110,
64'b1001100110011001011001100110011011000011001111001100001100111100,
64'b0000111111110000000011111111000001010101010101011010101010101010,
64'b0110100110010110011010011001011000110011110011000011001111001100,
64'b1010101010101010101010101010101010100101101001010101101001011010,
64'b1111000011110000111100001111000000000000000000000000000000000000,
64'b0110011010011001100110010110011011110000111100001111000011110000,
64'b1100110000110011001100111100110000110011110011000011001111001100,
64'b0000111100001111111100001111000011000011001111001100001100111100,
64'b0110100101101001100101101001011010100101010110101010010101011010,
64'b1010010110100101010110100101101000111100001111000011110000111100,
64'b1010010110100101010110100101101000000000111111111111111100000000,
64'b1100001100111100110000110011110011000011001111001100001100111100,
64'b0110100101101001100101101001011000111100001111000011110000111100,
64'b0101101001011010010110100101101011110000000011110000111111110000,
64'b0110100101101001100101101001011011001100110011001100110011001100,
64'b0110100110010110011010011001011010100101101001010101101001011010,
64'b1111111100000000111111110000000000110011110011000011001111001100,
64'b0101101010100101101001010101101010101010101010101010101010101010,
64'b1100001111000011001111000011110011111111000000001111111100000000,
64'b0101010101010101101010101010101000001111000011111111000011110000,
64'b0110011001100110011001100110011011110000000011110000111111110000,
64'b1010101010101010101010101010101011001100001100110011001111001100,
64'b0011110000111100001111000011110000001111111100000000111111110000,
64'b1010010101011010101001010101101011111111111111110000000000000000,
64'b0101101001011010010110100101101010100101010110101010010101011010,
64'b0110100110010110011010011001011010100101010110101010010101011010,
64'b1001100101100110100110010110011000000000111111111111111100000000,
64'b1100001100111100110000110011110001011010010110100101101001011010,
64'b1001011001101001011010011001011000110011110011000011001111001100,
64'b1111111111111111000000000000000010100101101001010101101001011010,
64'b1100110000110011001100111100110011001100110011001100110011001100,
64'b1010010101011010101001010101101011111111111111110000000000000000,
64'b0110011001100110011001100110011011111111000000001111111100000000,
64'b1001011010010110100101101001011010101010010101010101010110101010,
64'b1100110011001100110011001100110010100101101001010101101001011010,
64'b0000111111110000000011111111000010101010010101010101010110101010,
64'b1100110000110011001100111100110000000000000000000000000000000000,
64'b0011001111001100001100111100110010011001011001101001100101100110,
64'b0011110011000011110000110011110001100110100110011001100101100110,
64'b1100001111000011001111000011110011111111111111110000000000000000,
64'b1111000000001111000011111111000010011001011001101001100101100110,
64'b0011110011000011110000110011110000001111000011111111000011110000,
64'b1010101010101010101010101010101000110011110011000011001111001100,
64'b1010010110100101010110100101101001011010010110100101101001011010,
64'b0110011010011001100110010110011000000000000000000000000000000000,
64'b0011110000111100001111000011110001010101010101011010101010101010,
64'b1100001100111100110000110011110000110011001100111100110011001100,
64'b1111000011110000111100001111000010011001011001101001100101100110,
64'b0000000011111111111111110000000010011001100110010110011001100110,
64'b0000111100001111111100001111000010101010101010101010101010101010,
64'b0101101001011010010110100101101000111100001111000011110000111100,
64'b1111000000001111000011111111000001101001011010011001011010010110,
64'b1010010101011010101001010101101010101010101010101010101010101010,
64'b1010101001010101010101011010101001101001011010011001011010010110,
64'b0101101010100101101001010101101011111111000000001111111100000000,
64'b0110011001100110011001100110011010100101101001010101101001011010,
64'b0011001111001100001100111100110000110011110011000011001111001100,
64'b0110100101101001100101101001011000000000000000000000000000000000,
64'b1010010101011010101001010101101011001100110011001100110011001100,
64'b1111000000001111000011111111000001011010010110100101101001011010,
64'b1111111100000000111111110000000001101001011010011001011010010110,
64'b1111111111111111000000000000000000111100001111000011110000111100,
64'b0101010110101010010101011010101001100110011001100110011001100110,
64'b1001100101100110100110010110011000001111111100000000111111110000,
64'b0101101010100101101001010101101000000000111111111111111100000000,
64'b0011110000111100001111000011110011111111000000001111111100000000,
64'b1111000011110000111100001111000011111111111111110000000000000000,
64'b1111000000001111000011111111000011000011001111001100001100111100,
64'b0110100110010110011010011001011000111100001111000011110000111100,
64'b0101101010100101101001010101101001011010101001011010010101011010,
64'b1001011001101001011010011001011000000000000000000000000000000000,
64'b1111111111111111000000000000000011000011110000110011110000111100,
64'b1001100101100110100110010110011010011001100110010110011001100110,
64'b0011110011000011110000110011110011000011001111001100001100111100,
64'b0011110011000011110000110011110000001111000011111111000011110000,
64'b1001100101100110100110010110011010011001100110010110011001100110,
64'b1001100101100110100110010110011001010101101010100101010110101010,
64'b0011110000111100001111000011110001010101010101011010101010101010,
64'b1001100101100110100110010110011001010101010101011010101010101010,
64'b0000111111110000000011111111000000000000000000000000000000000000,
64'b1111000011110000111100001111000001011010101001011010010101011010,
64'b1111111111111111000000000000000000001111111100000000111111110000,
64'b1001011010010110100101101001011011001100001100110011001111001100,
64'b0000000000000000000000000000000010101010101010101010101010101010,
64'b0101010101010101101010101010101000001111111100000000111111110000,
64'b1111000000001111000011111111000010010110100101101001011010010110,
64'b1100110011001100110011001100110001011010101001011010010101011010,
64'b0110011001100110011001100110011011111111000000001111111100000000,
64'b1111000000001111000011111111000010010110100101101001011010010110,
64'b1010010101011010101001010101101001100110011001100110011001100110,
64'b1111111111111111000000000000000001100110011001100110011001100110,
64'b1111111111111111000000000000000001100110011001100110011001100110,
64'b1111000000001111000011111111000010101010101010101010101010101010,
64'b0000111100001111111100001111000011001100001100110011001111001100,
64'b0110100110010110011010011001011010101010010101010101010110101010,
64'b0011001100110011110011001100110000001111000011111111000011110000,
64'b1001011001101001011010011001011001100110011001100110011001100110,
64'b0011001100110011110011001100110000000000111111111111111100000000,
64'b0011001100110011110011001100110011000011001111001100001100111100,
64'b0110011010011001100110010110011011001100001100110011001111001100,
64'b0000000011111111111111110000000001010101010101011010101010101010,
64'b1001100110011001011001100110011011000011001111001100001100111100,
64'b0000000000000000000000000000000000111100001111000011110000111100,
64'b1010101010101010101010101010101010010110100101101001011010010110,
64'b1010101010101010101010101010101000111100001111000011110000111100,
64'b1010101001010101010101011010101011001100110011001100110011001100,
64'b0101010110101010010101011010101000001111000011111111000011110000,
64'b1001011001101001011010011001011010011001100110010110011001100110,
64'b1111000011110000111100001111000001010101101010100101010110101010,
64'b1001011001101001011010011001011010010110100101101001011010010110,
64'b0101101001011010010110100101101011111111111111110000000000000000,
64'b0101101001011010010110100101101001011010101001011010010101011010,
64'b0110100101101001100101101001011000001111000011111111000011110000,
64'b0101010101010101101010101010101001100110011001100110011001100110,
64'b1001011010010110100101101001011001011010101001011010010101011010,
64'b1010101010101010101010101010101000001111111100000000111111110000,
64'b1001011001101001011010011001011011000011001111001100001100111100,
64'b1111000011110000111100001111000000001111111100000000111111110000,
64'b1100001111000011001111000011110011110000111100001111000011110000,
64'b0110100110010110011010011001011011111111000000001111111100000000,
64'b0101010101010101101010101010101010010110100101101001011010010110,
64'b0000111100001111111100001111000010011001100110010110011001100110,
64'b1010101010101010101010101010101011000011001111001100001100111100,
64'b0110011010011001100110010110011000000000000000000000000000000000,
64'b1010101010101010101010101010101001100110100110011001100101100110,
64'b1111111111111111000000000000000001010101101010100101010110101010,
64'b0101101010100101101001010101101010010110100101101001011010010110,
64'b1111000011110000111100001111000011001100001100110011001111001100,
64'b0101010110101010010101011010101001010101101010100101010110101010,
64'b1100110011001100110011001100110001011010101001011010010101011010,
64'b0110100110010110011010011001011000000000111111111111111100000000,
64'b1111111100000000111111110000000011111111000000001111111100000000,
64'b0110011001100110011001100110011011111111111111110000000000000000,
64'b1010010101011010101001010101101011000011001111001100001100111100,
64'b0000111100001111111100001111000000111100001111000011110000111100,
64'b1111000000001111000011111111000001011010101001011010010101011010,
64'b0011110000111100001111000011110000000000000000000000000000000000,
64'b1111111100000000111111110000000011000011110000110011110000111100,
64'b0011110011000011110000110011110010011001100110010110011001100110,
64'b0101101001011010010110100101101011000011001111001100001100111100,
64'b1100110011001100110011001100110000001111000011111111000011110000,
64'b0101010110101010010101011010101001100110011001100110011001100110,
64'b0101101001011010010110100101101010010110100101101001011010010110,
64'b0011110011000011110000110011110001101001011010011001011010010110,
64'b1111111111111111000000000000000010100101101001010101101001011010,
64'b0011110000111100001111000011110011110000000011110000111111110000,
64'b1100110000110011001100111100110000110011001100111100110011001100,
64'b1111111100000000111111110000000001010101010101011010101010101010,
64'b1010101001010101010101011010101001011010010110100101101001011010,
64'b1010010101011010101001010101101001010101010101011010101010101010,
64'b1111111111111111000000000000000010010110100101101001011010010110,
64'b1111000000001111000011111111000010101010010101010101010110101010,
64'b1001100101100110100110010110011001100110011001100110011001100110,
64'b1111000011110000111100001111000001100110011001100110011001100110,
64'b1100110011001100110011001100110000001111111100000000111111110000,
64'b1100001111000011001111000011110010011001100110010110011001100110,
64'b1100110000110011001100111100110011111111000000001111111100000000,
64'b0101101001011010010110100101101001101001100101100110100110010110,
64'b0101010101010101101010101010101001011010010110100101101001011010,
64'b0110011010011001100110010110011000110011110011000011001111001100,
64'b0000111111110000000011111111000000111100110000111100001100111100,
64'b1010010101011010101001010101101000001111000011111111000011110000,
64'b1001100101100110100110010110011000110011001100111100110011001100,
64'b1001100101100110100110010110011011110000111100001111000011110000,
64'b1001011010010110100101101001011000001111111100000000111111110000,
64'b0101010110101010010101011010101010101010010101010101010110101010,
64'b0110011001100110011001100110011010100101010110101010010101011010,
64'b0110100110010110011010011001011001100110011001100110011001100110,
64'b1111111111111111000000000000000010010110100101101001011010010110,
64'b1001100110011001011001100110011001010101010101011010101010101010,
64'b0110100110010110011010011001011000111100110000111100001100111100,
64'b0011110011000011110000110011110000110011110011000011001111001100,
64'b0000000011111111111111110000000000001111000011111111000011110000,
64'b1111000011110000111100001111000011110000000011110000111111110000,
64'b0101101001011010010110100101101001010101101010100101010110101010,
64'b0011110000111100001111000011110001011010010110100101101001011010,
64'b0101101010100101101001010101101001010101101010100101010110101010,
64'b1111111111111111000000000000000000000000111111111111111100000000,
64'b0000111111110000000011111111000000110011001100111100110011001100,
64'b1010010101011010101001010101101001100110100110011001100101100110,
64'b0101101001011010010110100101101000111100001111000011110000111100,
64'b1010101010101010101010101010101001101001100101100110100110010110,
64'b1001011010010110100101101001011011001100110011001100110011001100,
64'b1001011001101001011010011001011001011010101001011010010101011010,
64'b1111000000001111000011111111000010100101101001010101101001011010,
64'b0101010101010101101010101010101011111111000000001111111100000000,
64'b0101010110101010010101011010101010101010010101010101010110101010,
64'b0011001111001100001100111100110010011001100110010110011001100110,
64'b0000111111110000000011111111000000110011110011000011001111001100,
64'b1100110000110011001100111100110000110011001100111100110011001100,
64'b1010101010101010101010101010101011111111111111110000000000000000,
64'b1010101001010101010101011010101001011010010110100101101001011010,
64'b1100110000110011001100111100110001101001011010011001011010010110,
64'b0011001111001100001100111100110010100101010110101010010101011010,
64'b0011110011000011110000110011110001100110011001100110011001100110,
64'b1111111100000000111111110000000011001100110011001100110011001100,
64'b1100110000110011001100111100110000111100110000111100001100111100,
64'b0101101001011010010110100101101001101001011010011001011010010110,
64'b0000111111110000000011111111000000111100110000111100001100111100,
64'b1100001100111100110000110011110001101001100101100110100110010110,
64'b1001100101100110100110010110011000000000111111111111111100000000,
64'b1111111100000000111111110000000001011010010110100101101001011010,
64'b1001011001101001011010011001011001101001100101100110100110010110,
64'b0101101010100101101001010101101010010110011010010110100110010110,
64'b0000111111110000000011111111000010100101101001010101101001011010,
64'b0011110011000011110000110011110001011010010110100101101001011010,
64'b1100001100111100110000110011110000000000000000000000000000000000,
64'b0000000000000000000000000000000000111100001111000011110000111100,
64'b0110100101101001100101101001011011110000111100001111000011110000,
64'b1111111111111111000000000000000011110000000011110000111111110000,
64'b0110100101101001100101101001011001101001100101100110100110010110,
64'b0110100101101001100101101001011001011010101001011010010101011010,
64'b1010101010101010101010101010101010010110011010010110100110010110,
64'b0101010110101010010101011010101011111111111111110000000000000000,
64'b0000000000000000000000000000000010011001011001101001100101100110,
64'b1010010110100101010110100101101000111100110000111100001100111100,
64'b0101101001011010010110100101101000111100110000111100001100111100,
64'b1001011010010110100101101001011010011001011001101001100101100110,
64'b0110100101101001100101101001011010011001011001101001100101100110,
64'b0011110000111100001111000011110000000000000000000000000000000000,
64'b1111000000001111000011111111000010100101010110101010010101011010,
64'b1111111100000000111111110000000011111111000000001111111100000000,
64'b0101101001011010010110100101101000000000111111111111111100000000,
64'b1001100110011001011001100110011010010110011010010110100110010110,
64'b0000000000000000000000000000000011001100001100110011001111001100,
64'b0011110011000011110000110011110010010110011010010110100110010110,
64'b1010010101011010101001010101101010101010101010101010101010101010,
64'b1111111111111111000000000000000001101001011010011001011010010110,
64'b1010101010101010101010101010101011110000000011110000111111110000,
64'b1010010110100101010110100101101001011010101001011010010101011010,
64'b1111111111111111000000000000000001101001011010011001011010010110,
64'b0101101001011010010110100101101011000011110000110011110000111100,
64'b0011110000111100001111000011110000000000000000000000000000000000,
64'b0000000011111111111111110000000001100110100110011001100101100110,
64'b0101010101010101101010101010101011111111111111110000000000000000,
64'b0011001111001100001100111100110011111111111111110000000000000000,
64'b0011110000111100001111000011110010010110011010010110100110010110,
64'b1010101010101010101010101010101010100101101001010101101001011010,
64'b1111000000001111000011111111000010010110011010010110100110010110,
64'b0110011010011001100110010110011001100110011001100110011001100110,
64'b0000000000000000000000000000000011000011001111001100001100111100,
64'b0110011001100110011001100110011010101010010101010101010110101010,
64'b0011001111001100001100111100110001100110100110011001100101100110,
64'b1010101010101010101010101010101001101001100101100110100110010110,
64'b1001100101100110100110010110011010100101010110101010010101011010,
64'b0000111111110000000011111111000010101010101010101010101010101010,
64'b0101010101010101101010101010101001101001011010011001011010010110,
64'b0110011001100110011001100110011010101010101010101010101010101010,
64'b1010010110100101010110100101101010101010101010101010101010101010,
64'b0000111111110000000011111111000010010110011010010110100110010110,
64'b1100110011001100110011001100110010011001011001101001100101100110,
64'b0000000011111111111111110000000010010110011010010110100110010110,
64'b0110100101101001100101101001011010010110100101101001011010010110,
64'b1010101010101010101010101010101011110000000011110000111111110000,
64'b0011110000111100001111000011110000110011001100111100110011001100,
64'b0000111100001111111100001111000001101001011010011001011010010110,
64'b1100110011001100110011001100110010010110011010010110100110010110,
64'b1100001111000011001111000011110011001100001100110011001111001100,
64'b1111111100000000111111110000000011001100110011001100110011001100,
64'b1100110011001100110011001100110011000011001111001100001100111100,
64'b1001011010010110100101101001011001100110011001100110011001100110,
64'b0011001111001100001100111100110011001100110011001100110011001100,
64'b1010101001010101010101011010101000111100110000111100001100111100,
64'b1111000011110000111100001111000001101001011010011001011010010110,
64'b1111111111111111000000000000000000111100110000111100001100111100,
64'b0110100110010110011010011001011001101001100101100110100110010110,
64'b0110011001100110011001100110011000000000111111111111111100000000,
64'b0000111111110000000011111111000001011010010110100101101001011010,
64'b1111111100000000111111110000000001101001100101100110100110010110,
64'b0101101001011010010110100101101010010110011010010110100110010110,
64'b0000111111110000000011111111000010100101101001010101101001011010,
64'b1010101010101010101010101010101001011010010110100101101001011010,
64'b0000000000000000000000000000000000111100001111000011110000111100,
64'b0011001100110011110011001100110010101010010101010101010110101010,
64'b1100110011001100110011001100110000111100110000111100001100111100,
64'b1001100110011001011001100110011010100101101001010101101001011010,
64'b1001011010010110100101101001011000110011001100111100110011001100,
64'b0000000011111111111111110000000000110011110011000011001111001100,
64'b1001011001101001011010011001011000001111000011111111000011110000,
64'b0011110011000011110000110011110011111111000000001111111100000000,
64'b0000000011111111111111110000000000000000111111111111111100000000,
64'b1111111100000000111111110000000000001111111100000000111111110000,
64'b0000111100001111111100001111000001011010101001011010010101011010,
64'b0000111100001111111100001111000010011001100110010110011001100110,
64'b1100001100111100110000110011110011001100110011001100110011001100,
64'b1010101010101010101010101010101010100101010110101010010101011010,
64'b1100001111000011001111000011110000110011001100111100110011001100,
64'b1001011010010110100101101001011001011010101001011010010101011010,
64'b1010010110100101010110100101101010011001011001101001100101100110,
64'b1111111100000000111111110000000001011010010110100101101001011010,
64'b1111111100000000111111110000000010100101101001010101101001011010,
64'b0000000000000000000000000000000011111111000000001111111100000000,
64'b0110011001100110011001100110011001010101010101011010101010101010,
64'b0101010110101010010101011010101011111111111111110000000000000000,
64'b1010101001010101010101011010101010101010010101010101010110101010,
64'b1111000000001111000011111111000011001100001100110011001111001100,
64'b0101101010100101101001010101101010010110100101101001011010010110,
64'b0110011001100110011001100110011001011010010110100101101001011010,
64'b0110011001100110011001100110011011001100001100110011001111001100,
64'b0011110011000011110000110011110011110000111100001111000011110000,
64'b1010010101011010101001010101101001100110100110011001100101100110,
64'b1010101001010101010101011010101001101001011010011001011010010110,
64'b1100001111000011001111000011110000110011110011000011001111001100,
64'b1111111100000000111111110000000000110011110011000011001111001100,
64'b1001011001101001011010011001011001010101010101011010101010101010,
64'b0000000011111111111111110000000011001100110011001100110011001100,
64'b0011001111001100001100111100110010101010101010101010101010101010,
64'b1100110000110011001100111100110010011001100110010110011001100110,
64'b1010010101011010101001010101101010100101101001010101101001011010,
64'b0110100110010110011010011001011001101001100101100110100110010110,
64'b0101010110101010010101011010101000110011110011000011001111001100,
64'b0011110000111100001111000011110000001111000011111111000011110000,
64'b1111000000001111000011111111000001010101101010100101010110101010,
64'b0110011010011001100110010110011011000011110000110011110000111100,
64'b0011001100110011110011001100110001101001100101100110100110010110,
64'b1010010101011010101001010101101010100101101001010101101001011010,
64'b0101010101010101101010101010101000001111000011111111000011110000,
64'b0011110011000011110000110011110011001100110011001100110011001100,
64'b0101010101010101101010101010101001011010010110100101101001011010,
64'b1010010110100101010110100101101011001100110011001100110011001100,
64'b0000111100001111111100001111000000111100001111000011110000111100,
64'b0110011010011001100110010110011010011001011001101001100101100110,
64'b0011110011000011110000110011110010010110011010010110100110010110,
64'b1100110011001100110011001100110011110000111100001111000011110000,
64'b0000111111110000000011111111000001010101101010100101010110101010,
64'b0011001111001100001100111100110010011001100110010110011001100110,
64'b1010010110100101010110100101101000001111111100000000111111110000,
64'b1100001111000011001111000011110010010110011010010110100110010110,
64'b1111000000001111000011111111000000110011110011000011001111001100,
64'b1100110000110011001100111100110001010101101010100101010110101010,
64'b1100110011001100110011001100110001011010010110100101101001011010,
64'b0101101010100101101001010101101000110011110011000011001111001100,
64'b1001100110011001011001100110011011110000111100001111000011110000,
64'b1010101010101010101010101010101000001111111100000000111111110000,
64'b0110011001100110011001100110011011000011110000110011110000111100,
64'b0101010110101010010101011010101000111100110000111100001100111100,
64'b1001100101100110100110010110011001010101101010100101010110101010,
64'b1010101001010101010101011010101010011001100110010110011001100110,
64'b0011110000111100001111000011110000111100001111000011110000111100,
64'b1111111100000000111111110000000010101010010101010101010110101010,
64'b0011110011000011110000110011110000111100110000111100001100111100,
64'b0011110011000011110000110011110010100101101001010101101001011010,
64'b1010010101011010101001010101101000110011001100111100110011001100,
64'b1100110000110011001100111100110000110011110011000011001111001100,
64'b1111000011110000111100001111000000001111000011111111000011110000,
64'b1001011001101001011010011001011011111111000000001111111100000000,
64'b1001100101100110100110010110011000000000111111111111111100000000,
64'b0011001100110011110011001100110000001111111100000000111111110000,
64'b0011110000111100001111000011110001011010101001011010010101011010,
64'b1111111100000000111111110000000001100110011001100110011001100110,
64'b1001100110011001011001100110011000111100001111000011110000111100,
64'b1010010101011010101001010101101010010110011010010110100110010110,
64'b1111111111111111000000000000000011111111111111110000000000000000,
64'b1111000000001111000011111111000011000011001111001100001100111100,
64'b0101101010100101101001010101101000001111111100000000111111110000,
64'b0110011010011001100110010110011001011010101001011010010101011010,
64'b0000111100001111111100001111000000110011110011000011001111001100,
64'b0101010110101010010101011010101011000011110000110011110000111100,
64'b0011110011000011110000110011110001010101101010100101010110101010,
64'b0110100101101001100101101001011000000000111111111111111100000000,
64'b1111000011110000111100001111000010100101010110101010010101011010,
64'b1010010101011010101001010101101011000011001111001100001100111100,
64'b0000000000000000000000000000000001010101101010100101010110101010,
64'b0011110000111100001111000011110010100101010110101010010101011010,
64'b0101010110101010010101011010101000001111111100000000111111110000,
64'b1100110011001100110011001100110001100110011001100110011001100110,
64'b0011001111001100001100111100110011000011001111001100001100111100,
64'b1111000000001111000011111111000010010110011010010110100110010110,
64'b0110100110010110011010011001011011001100110011001100110011001100,
64'b1100001111000011001111000011110000110011110011000011001111001100,
64'b1010010101011010101001010101101000110011001100111100110011001100,
64'b1111000011110000111100001111000010011001011001101001100101100110,
64'b1001011010010110100101101001011000000000111111111111111100000000,
64'b0101101010100101101001010101101001101001100101100110100110010110,
64'b1100001100111100110000110011110011111111000000001111111100000000,
64'b1100001100111100110000110011110000001111111100000000111111110000,
64'b1010010101011010101001010101101011001100001100110011001111001100,
64'b0000000000000000000000000000000000000000111111111111111100000000,
64'b0011110000111100001111000011110000111100001111000011110000111100,
64'b1001011010010110100101101001011011110000000011110000111111110000,
64'b1001011001101001011010011001011000111100110000111100001100111100,
64'b1001011010010110100101101001011001011010010110100101101001011010,
64'b1001100110011001011001100110011000001111000011111111000011110000,
64'b0101101001011010010110100101101011110000111100001111000011110000,
64'b1111111111111111000000000000000001101001011010011001011010010110,
64'b0011110000111100001111000011110011111111111111110000000000000000,
64'b1100001100111100110000110011110010010110011010010110100110010110,
64'b0101010110101010010101011010101011111111111111110000000000000000,
64'b1100110011001100110011001100110011111111000000001111111100000000,
64'b1100110000110011001100111100110000001111000011111111000011110000,
64'b0000000000000000000000000000000001010101010101011010101010101010,
64'b0000111111110000000011111111000010100101010110101010010101011010,
64'b1100001100111100110000110011110000000000111111111111111100000000,
64'b0011110011000011110000110011110001011010101001011010010101011010,
64'b0110100110010110011010011001011010011001011001101001100101100110,
64'b0011110000111100001111000011110011111111000000001111111100000000,
64'b1001100101100110100110010110011001010101101010100101010110101010,
64'b0000000000000000000000000000000011000011001111001100001100111100,
64'b1010010101011010101001010101101010101010101010101010101010101010,
64'b1111000000001111000011111111000010010110011010010110100110010110,
64'b0011001100110011110011001100110010101010101010101010101010101010,
64'b1111000011110000111100001111000010101010101010101010101010101010,
64'b1010010110100101010110100101101001010101101010100101010110101010,
64'b1001100110011001011001100110011001010101010101011010101010101010,
64'b1100110000110011001100111100110010101010010101010101010110101010,
64'b0110100110010110011010011001011001100110011001100110011001100110,
64'b0110011010011001100110010110011011110000000011110000111111110000,
64'b1001011010010110100101101001011001101001100101100110100110010110,
64'b1001100110011001011001100110011001101001100101100110100110010110,
64'b1111111100000000111111110000000000001111111100000000111111110000,
64'b0000000011111111111111110000000011110000111100001111000011110000,
64'b0011001100110011110011001100110000110011110011000011001111001100,
64'b0000111111110000000011111111000000110011110011000011001111001100,
64'b0101010101010101101010101010101001101001011010011001011010010110,
64'b1001011010010110100101101001011000001111111100000000111111110000,
64'b1001100101100110100110010110011000110011001100111100110011001100,
64'b1010010110100101010110100101101011001100110011001100110011001100,
64'b0110100101101001100101101001011010011001100110010110011001100110,
64'b0000111111110000000011111111000010010110100101101001011010010110,
64'b0101010101010101101010101010101000000000111111111111111100000000,
64'b0110100101101001100101101001011010010110011010010110100110010110,
64'b1010101001010101010101011010101000111100110000111100001100111100,
64'b0110100110010110011010011001011000000000111111111111111100000000,
64'b1111111100000000111111110000000011111111000000001111111100000000,
64'b1010010101011010101001010101101000001111000011111111000011110000,
64'b1010010101011010101001010101101000001111000011111111000011110000,
64'b1100001111000011001111000011110011000011001111001100001100111100,
64'b1010101010101010101010101010101001010101101010100101010110101010,
64'b1100001111000011001111000011110011110000111100001111000011110000,
64'b0000000011111111111111110000000001011010010110100101101001011010,
64'b1010010101011010101001010101101000111100001111000011110000111100,
64'b0011001111001100001100111100110001101001100101100110100110010110,
64'b0101101001011010010110100101101011111111111111110000000000000000,
64'b0110100101101001100101101001011010010110011010010110100110010110,
64'b0000111111110000000011111111000001011010101001011010010101011010,
64'b1010101010101010101010101010101001010101010101011010101010101010,
64'b1111111100000000111111110000000001010101010101011010101010101010,
64'b0011001100110011110011001100110011111111000000001111111100000000,
64'b1100001100111100110000110011110001010101101010100101010110101010,
64'b0000000011111111111111110000000001011010101001011010010101011010,
64'b1010010101011010101001010101101011001100110011001100110011001100,
64'b0000111111110000000011111111000011111111000000001111111100000000,
64'b0101010101010101101010101010101000110011110011000011001111001100,
64'b0110011010011001100110010110011000001111111100000000111111110000,
64'b0000111100001111111100001111000000111100110000111100001100111100,
64'b0011001111001100001100111100110000000000000000000000000000000000,
64'b1100001100111100110000110011110010010110011010010110100110010110,
64'b1010101001010101010101011010101001100110100110011001100101100110,
64'b1100110011001100110011001100110001100110011001100110011001100110,
64'b1111111111111111000000000000000001100110011001100110011001100110,
64'b1111000011110000111100001111000001010101010101011010101010101010,
64'b0101101010100101101001010101101000110011001100111100110011001100,
64'b1111111111111111000000000000000011001100001100110011001111001100,
64'b1001100101100110100110010110011001011010010110100101101001011010,
64'b1010101001010101010101011010101011111111111111110000000000000000,
64'b1100110011001100110011001100110000001111000011111111000011110000,
64'b0110100101101001100101101001011000000000111111111111111100000000,
64'b0101010110101010010101011010101011110000000011110000111111110000,
64'b1010010110100101010110100101101010101010101010101010101010101010,
64'b1111000000001111000011111111000000111100110000111100001100111100,
64'b0011001100110011110011001100110001101001011010011001011010010110,
64'b0101101001011010010110100101101010010110100101101001011010010110,
64'b0000000000000000000000000000000000111100001111000011110000111100,
64'b0101010110101010010101011010101011001100110011001100110011001100,
64'b1100110000110011001100111100110001011010010110100101101001011010,
64'b1010101010101010101010101010101010100101101001010101101001011010,
64'b1001011010010110100101101001011010011001011001101001100101100110,
64'b1001100110011001011001100110011000000000000000000000000000000000,
64'b0101101001011010010110100101101001010101101010100101010110101010,
64'b1100001100111100110000110011110001010101010101011010101010101010,
64'b1001100110011001011001100110011010101010010101010101010110101010,
64'b0011001111001100001100111100110001100110011001100110011001100110,
64'b1010101001010101010101011010101011110000000011110000111111110000,
64'b0101101001011010010110100101101001101001100101100110100110010110,
64'b1001100101100110100110010110011001101001100101100110100110010110,
64'b0000000000000000000000000000000000001111111100000000111111110000,
64'b0011001100110011110011001100110011110000111100001111000011110000,
64'b0000111100001111111100001111000000110011110011000011001111001100,
64'b0110011001100110011001100110011000110011110011000011001111001100,
64'b1100001100111100110000110011110010010110100101101001011010010110,
64'b0011001100110011110011001100110010010110011010010110100110010110,
64'b1010101001010101010101011010101011000011001111001100001100111100,
64'b0011001100110011110011001100110000111100001111000011110000111100,
64'b1100001100111100110000110011110001010101010101011010101010101010,
64'b0110011010011001100110010110011000110011110011000011001111001100,
64'b0110011001100110011001100110011000111100001111000011110000111100,
64'b0110011001100110011001100110011000110011110011000011001111001100,
64'b1010101010101010101010101010101011110000111100001111000011110000,
64'b1111000000001111000011111111000010101010010101010101010110101010,
64'b1010010101011010101001010101101001011010010110100101101001011010,
64'b0101010101010101101010101010101010011001011001101001100101100110,
64'b1001100101100110100110010110011010011001011001101001100101100110,
64'b0101101001011010010110100101101001101001100101100110100110010110,
64'b0110100101101001100101101001011000111100110000111100001100111100,
64'b0011001111001100001100111100110001011010101001011010010101011010,
64'b0110100101101001100101101001011000001111111100000000111111110000,
64'b1001100110011001011001100110011011001100110011001100110011001100,
64'b1010010101011010101001010101101010100101101001010101101001011010,
64'b1111000011110000111100001111000000001111111100000000111111110000,
64'b0101101001011010010110100101101000001111000011111111000011110000,
64'b0110011001100110011001100110011011111111000000001111111100000000,
64'b1111000011110000111100001111000000110011001100111100110011001100,
64'b1100001111000011001111000011110010011001011001101001100101100110,
64'b1001100110011001011001100110011011000011110000110011110000111100,
64'b1111000000001111000011111111000011000011110000110011110000111100,
64'b0110100110010110011010011001011011000011001111001100001100111100,
64'b1111000000001111000011111111000011110000000011110000111111110000,
64'b0000111111110000000011111111000001100110100110011001100101100110,
64'b1111000000001111000011111111000010101010010101010101010110101010,
64'b0101010110101010010101011010101011110000111100001111000011110000,
64'b0000000000000000000000000000000000110011110011000011001111001100,
64'b1001100101100110100110010110011010101010010101010101010110101010,
64'b0101010110101010010101011010101011111111000000001111111100000000,
64'b1001011010010110100101101001011001010101010101011010101010101010,
64'b0000111100001111111100001111000011110000111100001111000011110000,
64'b1010101010101010101010101010101001101001011010011001011010010110,
64'b1100001111000011001111000011110000001111111100000000111111110000,
64'b0011001100110011110011001100110010100101010110101010010101011010,
64'b0011001111001100001100111100110010100101010110101010010101011010,
64'b1010101001010101010101011010101010101010010101010101010110101010,
64'b1010101001010101010101011010101001101001011010011001011010010110,
64'b0000000011111111111111110000000010011001100110010110011001100110,
64'b1001100110011001011001100110011001010101101010100101010110101010,
64'b0000000000000000000000000000000000001111000011111111000011110000,
64'b1100001111000011001111000011110000110011001100111100110011001100,
64'b0011001100110011110011001100110001010101010101011010101010101010,
64'b1100001100111100110000110011110011001100110011001100110011001100,
64'b1111111100000000111111110000000001010101101010100101010110101010,
64'b0110011001100110011001100110011011000011001111001100001100111100,
64'b0000111111110000000011111111000010101010010101010101010110101010,
64'b0101101001011010010110100101101011001100001100110011001111001100,
64'b0101101001011010010110100101101000110011110011000011001111001100,
64'b0000000000000000000000000000000000110011001100111100110011001100,
64'b0011001111001100001100111100110001101001100101100110100110010110,
64'b0110011001100110011001100110011010010110100101101001011010010110,
64'b0101010110101010010101011010101010011001100110010110011001100110,
64'b1100110000110011001100111100110011111111000000001111111100000000,
64'b0110100110010110011010011001011001011010010110100101101001011010,
64'b0011110000111100001111000011110001100110011001100110011001100110,
64'b1111000000001111000011111111000001011010010110100101101001011010,
64'b0000111111110000000011111111000000110011001100111100110011001100,
64'b1001100101100110100110010110011011110000000011110000111111110000,
64'b0101010110101010010101011010101000110011001100111100110011001100,
64'b1010101010101010101010101010101010100101101001010101101001011010,
64'b0110100110010110011010011001011001011010010110100101101001011010,
64'b1001100110011001011001100110011001011010010110100101101001011010,
64'b1010010101011010101001010101101010010110011010010110100110010110,
64'b0000111100001111111100001111000011000011001111001100001100111100,
64'b1111000000001111000011111111000000111100001111000011110000111100,
64'b0110100110010110011010011001011001010101010101011010101010101010,
64'b1111000000001111000011111111000000110011110011000011001111001100,
64'b0110100110010110011010011001011000111100001111000011110000111100,
64'b1010101001010101010101011010101000110011110011000011001111001100,
64'b0101101001011010010110100101101011110000111100001111000011110000,
64'b0110011010011001100110010110011010101010010101010101010110101010,
64'b0110011001100110011001100110011001011010010110100101101001011010,
64'b0101010110101010010101011010101010011001011001101001100101100110,
64'b1001100101100110100110010110011010011001011001101001100101100110,
64'b1001011010010110100101101001011000000000111111111111111100000000,
64'b0110011010011001100110010110011010010110100101101001011010010110,
64'b1111111100000000111111110000000001101001100101100110100110010110,
64'b1010101001010101010101011010101011001100110011001100110011001100,
64'b1001011001101001011010011001011010101010010101010101010110101010,
64'b0000000011111111111111110000000011000011110000110011110000111100,
64'b1001011001101001011010011001011001101001100101100110100110010110,
64'b0011001100110011110011001100110010100101101001010101101001011010,
64'b1001100101100110100110010110011000001111000011111111000011110000,
64'b1100001111000011001111000011110010010110011010010110100110010110,
64'b1001011010010110100101101001011011001100001100110011001111001100,
64'b0011001100110011110011001100110001011010101001011010010101011010,
64'b0011110000111100001111000011110001100110011001100110011001100110,
64'b1111000000001111000011111111000001100110011001100110011001100110,
64'b0110100110010110011010011001011011000011110000110011110000111100,
64'b0110011001100110011001100110011000001111111100000000111111110000,
64'b1111000000001111000011111111000000110011110011000011001111001100,
64'b1111000011110000111100001111000001010101101010100101010110101010,
64'b0011001100110011110011001100110011000011001111001100001100111100,
64'b1111000000001111000011111111000011110000000011110000111111110000,
64'b1111000011110000111100001111000010011001011001101001100101100110,
64'b1001100101100110100110010110011010100101101001010101101001011010,
64'b1010101010101010101010101010101000110011001100111100110011001100,
64'b0011110011000011110000110011110011110000111100001111000011110000,
64'b0110100110010110011010011001011011111111111111110000000000000000,
64'b1111111100000000111111110000000011001100110011001100110011001100,
64'b1001100101100110100110010110011010010110100101101001011010010110,
64'b0011110000111100001111000011110000001111111100000000111111110000,
64'b0000111100001111111100001111000010101010010101010101010110101010,
64'b1100001111000011001111000011110000001111000011111111000011110000,
64'b0011001100110011110011001100110000110011001100111100110011001100,
64'b1001011010010110100101101001011011110000000011110000111111110000,
64'b1100110000110011001100111100110000000000111111111111111100000000,
64'b1111111100000000111111110000000001101001011010011001011010010110,
64'b0011001111001100001100111100110000110011110011000011001111001100,
64'b0110100110010110011010011001011001011010010110100101101001011010,
64'b1010010101011010101001010101101001010101101010100101010110101010,
64'b0000111100001111111100001111000000000000000000000000000000000000,
64'b0101101001011010010110100101101001011010010110100101101001011010,
64'b1100001111000011001111000011110001101001100101100110100110010110,
64'b0000111111110000000011111111000000000000111111111111111100000000,
64'b1111111100000000111111110000000000110011001100111100110011001100,
64'b1010010101011010101001010101101001010101101010100101010110101010,
64'b0101101001011010010110100101101001011010010110100101101001011010,
64'b0110100110010110011010011001011010101010010101010101010110101010,
64'b0000111100001111111100001111000001010101010101011010101010101010,
64'b0101010101010101101010101010101001101001100101100110100110010110,
64'b0000111100001111111100001111000010100101101001010101101001011010,
64'b0011110011000011110000110011110000110011110011000011001111001100,
64'b1100110000110011001100111100110000110011001100111100110011001100,
64'b1111111100000000111111110000000000000000000000000000000000000000,
64'b1001100101100110100110010110011000110011110011000011001111001100,
64'b0011110011000011110000110011110000001111111100000000111111110000,
64'b0000000000000000000000000000000001010101101010100101010110101010,
64'b1100110011001100110011001100110001101001011010011001011010010110,
64'b0000111100001111111100001111000001011010101001011010010101011010,
64'b0101010101010101101010101010101001010101010101011010101010101010,
64'b0101101010100101101001010101101001010101010101011010101010101010,
64'b1001100101100110100110010110011000000000000000000000000000000000,
64'b1100110011001100110011001100110000111100110000111100001100111100,
64'b1010010110100101010110100101101011000011110000110011110000111100,
64'b1111111111111111000000000000000000000000111111111111111100000000,
64'b1111000011110000111100001111000010100101101001010101101001011010,
64'b1100110000110011001100111100110000110011110011000011001111001100,
64'b0110011001100110011001100110011010101010101010101010101010101010,
64'b1100001100111100110000110011110010101010010101010101010110101010,
64'b0000000011111111111111110000000000110011001100111100110011001100,
64'b1100001111000011001111000011110011000011001111001100001100111100,
64'b0011110000111100001111000011110001100110100110011001100101100110,
64'b0000000011111111111111110000000001100110011001100110011001100110,
64'b0000000011111111111111110000000001100110011001100110011001100110,
64'b0000111100001111111100001111000010101010101010101010101010101010,
64'b0101101001011010010110100101101011110000000011110000111111110000,
64'b1100001111000011001111000011110010100101010110101010010101011010,
64'b0000111111110000000011111111000001010101010101011010101010101010,
64'b0000000011111111111111110000000010011001011001101001100101100110,
64'b1001011001101001011010011001011010100101101001010101101001011010,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b1100001100111100110000110011110010011001100110010110011001100110,
64'b0101010110101010010101011010101001011010010110100101101001011010,
64'b1001011001101001011010011001011001011010101001011010010101011010,
64'b0110011001100110011001100110011011000011110000110011110000111100,
64'b1001100101100110100110010110011010010110100101101001011010010110,
64'b0011001100110011110011001100110000111100001111000011110000111100,
64'b0011001111001100001100111100110011001100110011001100110011001100,
64'b0011001111001100001100111100110000000000111111111111111100000000,
64'b1111111111111111000000000000000001100110100110011001100101100110,
64'b0000111100001111111100001111000011001100110011001100110011001100,
64'b1010101010101010101010101010101001101001011010011001011010010110,
64'b0000111100001111111100001111000000110011110011000011001111001100,
64'b0000000000000000000000000000000001011010010110100101101001011010,
64'b0101101010100101101001010101101000111100001111000011110000111100,
64'b0011001100110011110011001100110010011001011001101001100101100110,
64'b0011110011000011110000110011110011001100001100110011001111001100,
64'b1001011010010110100101101001011010100101010110101010010101011010,
64'b1100001111000011001111000011110001101001100101100110100110010110,
64'b1111000011110000111100001111000000001111111100000000111111110000,
64'b1010010110100101010110100101101011110000111100001111000011110000,
64'b0000111100001111111100001111000011111111111111110000000000000000,
64'b0000000000000000000000000000000001101001011010011001011010010110,
64'b0101010110101010010101011010101001011010010110100101101001011010,
64'b0110011001100110011001100110011011000011001111001100001100111100,
64'b1111111100000000111111110000000010100101101001010101101001011010,
64'b1010101010101010101010101010101000110011110011000011001111001100,
64'b0110011010011001100110010110011000001111111100000000111111110000,
64'b0101101001011010010110100101101011000011110000110011110000111100,
64'b0101101010100101101001010101101000001111000011111111000011110000,
64'b0110100110010110011010011001011001100110100110011001100101100110,
64'b0000111111110000000011111111000000111100110000111100001100111100,
64'b0101010110101010010101011010101000000000111111111111111100000000,
64'b0011001111001100001100111100110011111111000000001111111100000000,
64'b0101010110101010010101011010101000000000000000000000000000000000,
64'b1010101010101010101010101010101001101001100101100110100110010110,
64'b0011001100110011110011001100110010011001011001101001100101100110,
64'b0011110000111100001111000011110011110000000011110000111111110000,
64'b1111111111111111000000000000000000110011110011000011001111001100,
64'b1100110011001100110011001100110001011010010110100101101001011010,
64'b1100001111000011001111000011110010101010010101010101010110101010,
64'b1001100101100110100110010110011000001111111100000000111111110000,
64'b1100110000110011001100111100110001010101101010100101010110101010,
64'b1001011001101001011010011001011001101001011010011001011010010110,
64'b0000000011111111111111110000000001011010101001011010010101011010,
64'b0011001100110011110011001100110001010101010101011010101010101010,
64'b0000111100001111111100001111000001010101010101011010101010101010,
64'b0011001100110011110011001100110000000000000000000000000000000000,
64'b1100110011001100110011001100110000111100110000111100001100111100,
64'b1111000011110000111100001111000011000011110000110011110000111100,
64'b1010010101011010101001010101101000000000111111111111111100000000,
64'b0000000000000000000000000000000010100101101001010101101001011010,
64'b0101101001011010010110100101101000110011110011000011001111001100,
64'b0101101001011010010110100101101010100101101001010101101001011010,
64'b0000000011111111111111110000000010010110100101101001011010010110,
64'b0011001111001100001100111100110000000000111111111111111100000000,
64'b0011001111001100001100111100110001101001011010011001011010010110,
64'b0000111100001111111100001111000011001100110011001100110011001100,
64'b0110100101101001100101101001011001010101010101011010101010101010,
64'b1100001100111100110000110011110000000000111111111111111100000000,
64'b1111000011110000111100001111000010101010010101010101010110101010,
64'b0110011001100110011001100110011010100101010110101010010101011010,
64'b1010101010101010101010101010101010011001100110010110011001100110,
64'b0110011001100110011001100110011001011010101001011010010101011010,
64'b0000111111110000000011111111000000110011001100111100110011001100,
64'b0000111111110000000011111111000000111100001111000011110000111100,
64'b0110100110010110011010011001011010011001011001101001100101100110,
64'b1111111100000000111111110000000001101001100101100110100110010110,
64'b1001011001101001011010011001011011111111111111110000000000000000,
64'b0011110011000011110000110011110001101001100101100110100110010110,
64'b1111000000001111000011111111000001011010010110100101101001011010,
64'b0000000011111111111111110000000011001100110011001100110011001100,
64'b1001100110011001011001100110011001010101010101011010101010101010,
64'b0000111111110000000011111111000010011001100110010110011001100110,
64'b0101101001011010010110100101101001100110100110011001100101100110,
64'b0110011001100110011001100110011000111100001111000011110000111100,
64'b0101101001011010010110100101101001100110100110011001100101100110,
64'b0000111100001111111100001111000001011010010110100101101001011010,
64'b1111000011110000111100001111000010100101010110101010010101011010,
64'b1100110000110011001100111100110001101001011010011001011010010110,
64'b1111111100000000111111110000000000111100110000111100001100111100,
64'b0000111100001111111100001111000000000000000000000000000000000000,
64'b0110100101101001100101101001011010010110011010010110100110010110,
64'b1010010101011010101001010101101000110011110011000011001111001100,
64'b0011110000111100001111000011110011110000111100001111000011110000,
64'b0101010110101010010101011010101011001100110011001100110011001100,
64'b0101101010100101101001010101101010010110100101101001011010010110,
64'b0101010110101010010101011010101001101001011010011001011010010110,
64'b1001011010010110100101101001011010100101010110101010010101011010,
64'b0101010110101010010101011010101011000011110000110011110000111100,
64'b1111000011110000111100001111000010011001011001101001100101100110,
64'b0101101001011010010110100101101000110011110011000011001111001100,
64'b1010010110100101010110100101101001101001100101100110100110010110,
64'b0101010101010101101010101010101001011010101001011010010101011010,
64'b1111111100000000111111110000000010101010101010101010101010101010,
64'b0110100110010110011010011001011000111100110000111100001100111100,
64'b0110011010011001100110010110011010100101101001010101101001011010,
64'b0000111111110000000011111111000011111111000000001111111100000000,
64'b0011001100110011110011001100110011110000111100001111000011110000,
64'b1100110000110011001100111100110011000011001111001100001100111100,
64'b1001100110011001011001100110011011000011001111001100001100111100,
64'b1100001100111100110000110011110001100110100110011001100101100110,
64'b0011001100110011110011001100110000001111111100000000111111110000,
64'b1111111100000000111111110000000001101001011010011001011010010110,
64'b0011001111001100001100111100110011110000111100001111000011110000,
64'b0110100110010110011010011001011010010110011010010110100110010110,
64'b0110011010011001100110010110011011001100001100110011001111001100,
64'b0110011010011001100110010110011001100110011001100110011001100110,
64'b0000111100001111111100001111000011110000000011110000111111110000,
64'b1100110011001100110011001100110010011001011001101001100101100110,
64'b1100001100111100110000110011110001010101010101011010101010101010,
64'b0011001111001100001100111100110011111111000000001111111100000000,
64'b0101010101010101101010101010101011110000000011110000111111110000,
64'b1111000011110000111100001111000011110000000011110000111111110000,
64'b1111000000001111000011111111000011000011110000110011110000111100,
64'b1001011010010110100101101001011010101010010101010101010110101010,
64'b0101101010100101101001010101101011000011001111001100001100111100,
64'b1111111100000000111111110000000001010101101010100101010110101010,
64'b1100110000110011001100111100110000111100110000111100001100111100,
64'b1100001100111100110000110011110010100101101001010101101001011010,
64'b0101101010100101101001010101101010010110100101101001011010010110,
64'b0110011001100110011001100110011000000000111111111111111100000000,
64'b0101010101010101101010101010101001101001011010011001011010010110,
64'b1001100101100110100110010110011011001100110011001100110011001100,
64'b1100110000110011001100111100110001010101010101011010101010101010,
64'b0011110000111100001111000011110000000000111111111111111100000000,
64'b0011001111001100001100111100110010101010010101010101010110101010,
64'b1010101001010101010101011010101010100101010110101010010101011010,
64'b0000111111110000000011111111000010011001100110010110011001100110,
64'b1100001111000011001111000011110001011010101001011010010101011010,
64'b1010010101011010101001010101101011001100110011001100110011001100,
64'b1010010110100101010110100101101000000000111111111111111100000000,
64'b0101101010100101101001010101101010011001100110010110011001100110,
64'b1100110000110011001100111100110001011010010110100101101001011010,
64'b1001011010010110100101101001011011001100001100110011001111001100,
64'b1100110011001100110011001100110001100110100110011001100101100110,
64'b0110100101101001100101101001011000110011001100111100110011001100,
64'b0000111100001111111100001111000000001111111100000000111111110000,
64'b1010010101011010101001010101101010100101101001010101101001011010,
64'b0000111100001111111100001111000011111111111111110000000000000000,
64'b0011001100110011110011001100110011001100001100110011001111001100,
64'b1010101001010101010101011010101001011010010110100101101001011010,
64'b0000111111110000000011111111000001101001011010011001011010010110,
64'b1001100101100110100110010110011001010101101010100101010110101010,
64'b0110100110010110011010011001011010100101101001010101101001011010,
64'b0110011001100110011001100110011010010110011010010110100110010110,
64'b1001011001101001011010011001011010101010101010101010101010101010,
64'b0101101001011010010110100101101000111100110000111100001100111100,
64'b1111111111111111000000000000000001100110011001100110011001100110,
64'b1010101001010101010101011010101000110011001100111100110011001100,
64'b1001011010010110100101101001011001101001011010011001011010010110,
64'b1001011001101001011010011001011011000011001111001100001100111100,
64'b1001100101100110100110010110011011001100110011001100110011001100,
64'b1111000011110000111100001111000000001111000011111111000011110000,
64'b1111111111111111000000000000000011111111000000001111111100000000,
64'b1010010110100101010110100101101011001100110011001100110011001100,
64'b0011001111001100001100111100110001101001100101100110100110010110,
64'b1100110000110011001100111100110000110011110011000011001111001100,
64'b0011110011000011110000110011110010010110011010010110100110010110,
64'b0000111100001111111100001111000001100110011001100110011001100110,
64'b1010101010101010101010101010101011110000000011110000111111110000,
64'b0000111100001111111100001111000010010110100101101001011010010110,
64'b1111000011110000111100001111000011110000111100001111000011110000,
64'b1010101010101010101010101010101001101001100101100110100110010110,
64'b1100110000110011001100111100110001011010101001011010010101011010,
64'b0000111100001111111100001111000011110000111100001111000011110000,
64'b0101010110101010010101011010101011111111000000001111111100000000,
64'b0110011001100110011001100110011001010101010101011010101010101010,
64'b1001011010010110100101101001011011110000111100001111000011110000,
64'b0101010110101010010101011010101011000011001111001100001100111100,
64'b0000111100001111111100001111000000001111000011111111000011110000,
64'b0101101010100101101001010101101000111100110000111100001100111100,
64'b0101010110101010010101011010101010010110100101101001011010010110,
64'b0110011001100110011001100110011000000000111111111111111100000000,
64'b1111111100000000111111110000000001101001100101100110100110010110,
64'b0101010110101010010101011010101011111111000000001111111100000000,
64'b1100110011001100110011001100110000111100110000111100001100111100,
64'b0000111100001111111100001111000011001100001100110011001111001100,
64'b0101010110101010010101011010101001010101101010100101010110101010,
64'b1001100110011001011001100110011011111111111111110000000000000000,
64'b0011110000111100001111000011110011001100110011001100110011001100,
64'b1100001100111100110000110011110001010101101010100101010110101010,
64'b1100110011001100110011001100110000001111111100000000111111110000,
64'b0000111111110000000011111111000000001111111100000000111111110000,
64'b0110011001100110011001100110011001011010010110100101101001011010,
64'b1010101001010101010101011010101001011010010110100101101001011010,
64'b0000111111110000000011111111000011001100001100110011001111001100,
64'b1111000011110000111100001111000010011001011001101001100101100110,
64'b0101101001011010010110100101101010010110100101101001011010010110,
64'b0011001111001100001100111100110000110011001100111100110011001100,
64'b0000111111110000000011111111000001010101010101011010101010101010,
64'b1111111111111111000000000000000011111111111111110000000000000000,
64'b1001011010010110100101101001011010101010101010101010101010101010,
64'b1100001100111100110000110011110000111100001111000011110000111100,
64'b1111111111111111000000000000000000111100110000111100001100111100,
64'b1111111100000000111111110000000011110000111100001111000011110000,
64'b0101101010100101101001010101101000000000111111111111111100000000,
64'b0011110011000011110000110011110000110011110011000011001111001100,
64'b0000000011111111111111110000000000110011110011000011001111001100,
64'b1001100110011001011001100110011000001111000011111111000011110000,
64'b1111000000001111000011111111000001101001011010011001011010010110,
64'b0101101010100101101001010101101011000011001111001100001100111100,
64'b1100110000110011001100111100110011110000111100001111000011110000,
64'b1111000000001111000011111111000001100110011001100110011001100110,
64'b0110011001100110011001100110011010101010101010101010101010101010,
64'b1100001100111100110000110011110001100110011001100110011001100110,
64'b1001011001101001011010011001011000001111111100000000111111110000,
64'b0000111111110000000011111111000011110000000011110000111111110000,
64'b1010010101011010101001010101101001010101101010100101010110101010,
64'b1001011001101001011010011001011011111111111111110000000000000000,
64'b0101101001011010010110100101101010100101101001010101101001011010,
64'b0110011010011001100110010110011000001111000011111111000011110000,
64'b1010010101011010101001010101101011111111000000001111111100000000,
64'b1010010101011010101001010101101001101001100101100110100110010110,
64'b0000111111110000000011111111000001011010101001011010010101011010,
64'b0110011010011001100110010110011011111111000000001111111100000000,
64'b0101101010100101101001010101101000111100001111000011110000111100,
64'b1111000011110000111100001111000011001100110011001100110011001100,
64'b0101101010100101101001010101101000111100001111000011110000111100,
64'b0101101010100101101001010101101000000000111111111111111100000000,
64'b1010010110100101010110100101101000000000111111111111111100000000,
64'b0011110000111100001111000011110001100110011001100110011001100110,
64'b0011110011000011110000110011110000000000000000000000000000000000,
64'b1001100101100110100110010110011010011001011001101001100101100110,
64'b1100001111000011001111000011110001010101101010100101010110101010,
64'b0110011010011001100110010110011001010101010101011010101010101010,
64'b1100110000110011001100111100110000111100110000111100001100111100,
64'b0000000011111111111111110000000011001100001100110011001111001100,
64'b1100001111000011001111000011110001010101010101011010101010101010,
64'b0110011010011001100110010110011000001111111100000000111111110000,
64'b0101010110101010010101011010101011110000111100001111000011110000,
64'b1100110000110011001100111100110000001111111100000000111111110000,
64'b0110011010011001100110010110011011111111111111110000000000000000,
64'b1001100101100110100110010110011001010101010101011010101010101010,
64'b1010010101011010101001010101101010010110100101101001011010010110,
64'b1111000000001111000011111111000010101010101010101010101010101010,
64'b0110100101101001100101101001011011000011110000110011110000111100,
64'b0000111111110000000011111111000000110011001100111100110011001100,
64'b0110100101101001100101101001011011001100110011001100110011001100,
64'b1010010110100101010110100101101001011010101001011010010101011010,
64'b0101010101010101101010101010101010100101101001010101101001011010,
64'b1010010101011010101001010101101001100110011001100110011001100110,
64'b0110100101101001100101101001011010101010010101010101010110101010,
64'b1001100110011001011001100110011011111111000000001111111100000000,
64'b0000111100001111111100001111000000000000111111111111111100000000,
64'b0110100101101001100101101001011000000000000000000000000000000000,
64'b0110100101101001100101101001011001100110011001100110011001100110,
64'b0011001111001100001100111100110001101001100101100110100110010110,
64'b0000000011111111111111110000000011001100110011001100110011001100,
64'b0110100110010110011010011001011000001111111100000000111111110000,
64'b1010101001010101010101011010101001011010010110100101101001011010,
64'b1100001100111100110000110011110001011010010110100101101001011010,
64'b1001100101100110100110010110011011001100001100110011001111001100,
64'b0110011001100110011001100110011010011001011001101001100101100110,
64'b0110011010011001100110010110011010010110100101101001011010010110,
64'b1100001100111100110000110011110000110011001100111100110011001100,
64'b1001011010010110100101101001011001010101010101011010101010101010,
64'b0101010110101010010101011010101011111111111111110000000000000000,
64'b0110100110010110011010011001011010101010101010101010101010101010,
64'b0110100110010110011010011001011000111100001111000011110000111100,
64'b0101101001011010010110100101101011000011001111001100001100111100,
64'b1001100110011001011001100110011010100101101001010101101001011010,
64'b1111111100000000111111110000000010101010101010101010101010101010,
64'b0101010101010101101010101010101000001111111100000000111111110000,
64'b0000111100001111111100001111000010010110011010010110100110010110,
64'b1001100110011001011001100110011000110011001100111100110011001100,
64'b0101010101010101101010101010101001100110100110011001100101100110,
64'b0110100101101001100101101001011000111100001111000011110000111100,
64'b0110011001100110011001100110011000001111111100000000111111110000,
64'b1111000000001111000011111111000011110000111100001111000011110000,
64'b0110100101101001100101101001011000111100001111000011110000111100,
64'b1010010110100101010110100101101011001100001100110011001111001100,
64'b0110100110010110011010011001011001101001011010011001011010010110,
64'b0000111111110000000011111111000011001100110011001100110011001100,
64'b0000111100001111111100001111000000110011110011000011001111001100,
64'b1010101001010101010101011010101001100110011001100110011001100110,
64'b1001100110011001011001100110011000000000111111111111111100000000,
64'b0101101010100101101001010101101000111100110000111100001100111100,
64'b0000111100001111111100001111000001011010010110100101101001011010,
64'b0011001100110011110011001100110001101001011010011001011010010110,
64'b0000000011111111111111110000000010100101010110101010010101011010,
64'b1111000011110000111100001111000000000000111111111111111100000000,
64'b1111000011110000111100001111000011111111000000001111111100000000,
64'b0000000011111111111111110000000000001111111100000000111111110000,
64'b0011110011000011110000110011110000001111000011111111000011110000,
64'b1111111111111111000000000000000001101001100101100110100110010110,
64'b1111000011110000111100001111000001011010010110100101101001011010,
64'b0110011010011001100110010110011010100101101001010101101001011010,
64'b0110011010011001100110010110011000111100001111000011110000111100,
64'b1100001111000011001111000011110011111111111111110000000000000000,
64'b0110100110010110011010011001011001011010101001011010010101011010,
64'b1100110000110011001100111100110010011001011001101001100101100110,
64'b0000111100001111111100001111000011000011001111001100001100111100,
64'b0011110000111100001111000011110001100110100110011001100101100110,
64'b0011001111001100001100111100110011111111111111110000000000000000,
64'b0000111100001111111100001111000001010101010101011010101010101010,
64'b1001011010010110100101101001011000000000111111111111111100000000,
64'b1111111100000000111111110000000011111111000000001111111100000000,
64'b1100001100111100110000110011110010010110011010010110100110010110,
64'b0101101001011010010110100101101000110011110011000011001111001100,
64'b1100001111000011001111000011110010011001011001101001100101100110,
64'b0110100101101001100101101001011010100101010110101010010101011010,
64'b1010010101011010101001010101101000000000000000000000000000000000,
64'b1001011001101001011010011001011001100110100110011001100101100110,
64'b0000111100001111111100001111000001101001011010011001011010010110,
64'b0101010110101010010101011010101011110000000011110000111111110000,
64'b1010010101011010101001010101101011000011110000110011110000111100,
64'b0000111100001111111100001111000010101010101010101010101010101010,
64'b1111111100000000111111110000000001100110011001100110011001100110,
64'b0110100110010110011010011001011001010101010101011010101010101010,
64'b1111111111111111000000000000000001010101010101011010101010101010,
64'b1111000000001111000011111111000000111100110000111100001100111100,
64'b0011001111001100001100111100110001011010010110100101101001011010,
64'b0011110011000011110000110011110011000011110000110011110000111100,
64'b1001011010010110100101101001011011001100001100110011001111001100,
64'b0011001111001100001100111100110000000000000000000000000000000000,
64'b0011001111001100001100111100110011000011110000110011110000111100,
64'b1100110000110011001100111100110001101001100101100110100110010110,
64'b1100110011001100110011001100110010101010010101010101010110101010,
64'b1010010101011010101001010101101010100101010110101010010101011010,
64'b1001100101100110100110010110011001100110011001100110011001100110,
64'b1010010101011010101001010101101000111100001111000011110000111100,
64'b0101010110101010010101011010101011001100110011001100110011001100,
64'b1010010110100101010110100101101001100110011001100110011001100110,
64'b1100001111000011001111000011110001011010101001011010010101011010,
64'b0101010110101010010101011010101010011001011001101001100101100110,
64'b1100001100111100110000110011110010100101010110101010010101011010,
64'b1001011010010110100101101001011010100101101001010101101001011010,
64'b0101101001011010010110100101101010101010101010101010101010101010,
64'b0000000000000000000000000000000000001111111100000000111111110000,
64'b1001011010010110100101101001011010010110011010010110100110010110,
64'b0000111100001111111100001111000000110011001100111100110011001100,
64'b1010010101011010101001010101101001100110100110011001100101100110,
64'b1010010110100101010110100101101000111100001111000011110000111100,
64'b0011110000111100001111000011110000001111111100000000111111110000,
64'b0101101001011010010110100101101011110000111100001111000011110000,
64'b1001011001101001011010011001011000111100001111000011110000111100,
64'b1100110011001100110011001100110011001100001100110011001111001100,
64'b0110100110010110011010011001011010010110100101101001011010010110,
64'b0101101010100101101001010101101001010101101010100101010110101010,
64'b1100001100111100110000110011110011001100110011001100110011001100,
64'b0011001111001100001100111100110000110011001100111100110011001100,
64'b0000000000000000000000000000000000001111111100000000111111110000,
64'b1100001100111100110000110011110010100101010110101010010101011010,
64'b1111111100000000111111110000000000001111000011111111000011110000,
64'b0110011010011001100110010110011000000000000000000000000000000000,
64'b0011001111001100001100111100110011000011001111001100001100111100,
64'b1010010101011010101001010101101011110000111100001111000011110000,
64'b0011001111001100001100111100110010010110011010010110100110010110,
64'b0011110011000011110000110011110010101010010101010101010110101010,
64'b0101101001011010010110100101101001100110100110011001100101100110,
64'b1100001100111100110000110011110001100110011001100110011001100110,
64'b1111111100000000111111110000000000000000000000000000000000000000,
64'b1010010110100101010110100101101000001111111100000000111111110000,
64'b0101101001011010010110100101101010100101101001010101101001011010,
64'b0000111100001111111100001111000010100101010110101010010101011010,
64'b0110100110010110011010011001011001010101101010100101010110101010,
64'b1010101010101010101010101010101010101010010101010101010110101010,
64'b1010101010101010101010101010101011000011110000110011110000111100,
64'b1100001111000011001111000011110010010110011010010110100110010110,
64'b0011110000111100001111000011110000001111000011111111000011110000,
64'b0110011001100110011001100110011001010101101010100101010110101010,
64'b0101010110101010010101011010101000111100001111000011110000111100,
64'b1111000011110000111100001111000000000000111111111111111100000000,
64'b0000000000000000000000000000000010011001011001101001100101100110,
64'b1100110011001100110011001100110010101010101010101010101010101010,
64'b1100110011001100110011001100110000000000111111111111111100000000,
64'b1100110000110011001100111100110000110011110011000011001111001100,
64'b1111000000001111000011111111000001100110100110011001100101100110,
64'b0000111111110000000011111111000000110011001100111100110011001100,
64'b1001100110011001011001100110011000110011001100111100110011001100,
64'b1010010110100101010110100101101010100101010110101010010101011010,
64'b0110100110010110011010011001011010010110011010010110100110010110,
64'b0101010101010101101010101010101001010101101010100101010110101010,
64'b0101010101010101101010101010101010011001100110010110011001100110,
64'b1001011010010110100101101001011000001111111100000000111111110000,
64'b1001011010010110100101101001011011111111111111110000000000000000,
64'b0000111111110000000011111111000010010110100101101001011010010110,
64'b0101101001011010010110100101101001100110011001100110011001100110,
64'b1111000011110000111100001111000011111111111111110000000000000000,
64'b0000111100001111111100001111000010100101101001010101101001011010,
64'b1010101001010101010101011010101011000011110000110011110000111100,
64'b1010101001010101010101011010101001011010010110100101101001011010,
64'b0011110000111100001111000011110001011010010110100101101001011010,
64'b1001100101100110100110010110011001100110100110011001100101100110,
64'b1001011001101001011010011001011000111100110000111100001100111100,
64'b1100110011001100110011001100110010011001100110010110011001100110,
64'b0110011001100110011001100110011000111100001111000011110000111100,
64'b0110100110010110011010011001011010101010010101010101010110101010,
64'b1100001100111100110000110011110000000000000000000000000000000000,
64'b1111111100000000111111110000000001101001100101100110100110010110,
64'b1010101001010101010101011010101000001111000011111111000011110000,
64'b0000000000000000000000000000000011111111000000001111111100000000,
64'b1010101001010101010101011010101011001100001100110011001111001100,
64'b1001011010010110100101101001011010101010010101010101010110101010,
64'b0000000000000000000000000000000000000000111111111111111100000000,
64'b1111000000001111000011111111000001100110100110011001100101100110,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b0101101010100101101001010101101000111100110000111100001100111100,
64'b1010101001010101010101011010101001100110100110011001100101100110,
64'b0101010101010101101010101010101011001100001100110011001111001100,
64'b1001100101100110100110010110011010010110100101101001011010010110,
64'b1001100110011001011001100110011011000011001111001100001100111100,
64'b0000111111110000000011111111000011001100110011001100110011001100,
64'b0000000000000000000000000000000011111111000000001111111100000000,
64'b0101010110101010010101011010101001010101010101011010101010101010,
64'b0110011001100110011001100110011000001111000011111111000011110000,
64'b0110011010011001100110010110011010011001100110010110011001100110,
64'b1001100110011001011001100110011001010101010101011010101010101010,
64'b0101010110101010010101011010101001101001011010011001011010010110,
64'b0000111100001111111100001111000001100110011001100110011001100110,
64'b1010101001010101010101011010101011110000000011110000111111110000,
64'b0110100110010110011010011001011001101001011010011001011010010110,
64'b0000111100001111111100001111000010100101101001010101101001011010,
64'b1100110011001100110011001100110001101001100101100110100110010110,
64'b0101010110101010010101011010101011110000000011110000111111110000,
64'b0101101001011010010110100101101011110000111100001111000011110000,
64'b0011001100110011110011001100110001010101010101011010101010101010,
64'b1100110000110011001100111100110011001100110011001100110011001100,
64'b0110100101101001100101101001011001010101101010100101010110101010,
64'b1100110011001100110011001100110010010110100101101001011010010110,
64'b0000111100001111111100001111000001100110011001100110011001100110,
64'b1100110011001100110011001100110001101001100101100110100110010110,
64'b1001011001101001011010011001011010010110100101101001011010010110,
64'b1111111111111111000000000000000000000000111111111111111100000000,
64'b0110011001100110011001100110011001101001100101100110100110010110,
64'b1001011001101001011010011001011010011001011001101001100101100110,
64'b1111111111111111000000000000000010010110011010010110100110010110,
64'b0101101010100101101001010101101000000000111111111111111100000000,
64'b0011110000111100001111000011110001010101101010100101010110101010,
64'b1111000011110000111100001111000011001100110011001100110011001100,
64'b1010010110100101010110100101101001011010010110100101101001011010,
64'b0110100110010110011010011001011000110011001100111100110011001100,
64'b0101101001011010010110100101101011000011001111001100001100111100,
64'b1111111100000000111111110000000000111100001111000011110000111100,
64'b0101101001011010010110100101101000111100110000111100001100111100,
64'b0011110011000011110000110011110011000011001111001100001100111100,
64'b1010101010101010101010101010101011111111111111110000000000000000,
64'b1001011010010110100101101001011010010110011010010110100110010110,
64'b0011110011000011110000110011110011000011110000110011110000111100,
64'b1010101010101010101010101010101000111100110000111100001100111100,
64'b0110011010011001100110010110011001010101010101011010101010101010,
64'b1010010101011010101001010101101001100110011001100110011001100110,
64'b0101010110101010010101011010101011110000111100001111000011110000,
64'b0011001111001100001100111100110000110011110011000011001111001100,
64'b1001011001101001011010011001011011110000111100001111000011110000,
64'b0011001111001100001100111100110001011010101001011010010101011010,
64'b1111111111111111000000000000000000001111111100000000111111110000,
64'b0011001111001100001100111100110011110000000011110000111111110000,
64'b1111000000001111000011111111000001011010101001011010010101011010,
64'b0110011001100110011001100110011000000000000000000000000000000000,
64'b1100001100111100110000110011110010010110011010010110100110010110,
64'b1111000000001111000011111111000010100101010110101010010101011010,
64'b0110011001100110011001100110011001011010101001011010010101011010,
64'b1100001111000011001111000011110001100110011001100110011001100110,
64'b1001100101100110100110010110011010010110100101101001011010010110,
64'b1001100110011001011001100110011001010101101010100101010110101010,
64'b0000111100001111111100001111000000001111000011111111000011110000,
64'b0011110011000011110000110011110011111111000000001111111100000000,
64'b1010010110100101010110100101101011001100001100110011001111001100,
64'b0000000000000000000000000000000010101010010101010101010110101010,
64'b1010010110100101010110100101101000000000111111111111111100000000,
64'b0000000011111111111111110000000001100110100110011001100101100110,
64'b1001011010010110100101101001011010101010101010101010101010101010,
64'b1111000000001111000011111111000000111100110000111100001100111100,
64'b0000000011111111111111110000000001100110100110011001100101100110,
64'b1001011010010110100101101001011011001100001100110011001111001100,
64'b0000111111110000000011111111000010010110100101101001011010010110,
64'b1001011010010110100101101001011011000011001111001100001100111100,
64'b0101010110101010010101011010101010010110011010010110100110010110,
64'b1111111100000000111111110000000000000000111111111111111100000000,
64'b0110100101101001100101101001011011110000000011110000111111110000,
64'b0000111111110000000011111111000010010110011010010110100110010110,
64'b0000111100001111111100001111000011000011110000110011110000111100,
64'b0110011010011001100110010110011010101010101010101010101010101010,
64'b0011110000111100001111000011110000110011110011000011001111001100,
64'b1100001111000011001111000011110011001100001100110011001111001100,
64'b0011001111001100001100111100110000111100110000111100001100111100,
64'b1111000000001111000011111111000011110000111100001111000011110000,
64'b0110011001100110011001100110011011111111111111110000000000000000,
64'b0000000011111111111111110000000001101001100101100110100110010110,
64'b1001100101100110100110010110011000001111111100000000111111110000,
64'b1100110000110011001100111100110000111100110000111100001100111100,
64'b0000000011111111111111110000000001010101010101011010101010101010,
64'b1010101001010101010101011010101010101010010101010101010110101010,
64'b1010010110100101010110100101101010010110011010010110100110010110,
64'b1111000000001111000011111111000010100101010110101010010101011010,
64'b0000111111110000000011111111000001100110011001100110011001100110,
64'b1001100101100110100110010110011000001111000011111111000011110000,
64'b1100110000110011001100111100110000001111000011111111000011110000,
64'b1001011001101001011010011001011001011010101001011010010101011010,
64'b1111000011110000111100001111000001010101101010100101010110101010,
64'b1111000011110000111100001111000000000000000000000000000000000000,
64'b1111111100000000111111110000000010010110011010010110100110010110,
64'b0000111111110000000011111111000011111111000000001111111100000000,
64'b0101101010100101101001010101101011110000000011110000111111110000,
64'b1010101001010101010101011010101001100110011001100110011001100110,
64'b1111000011110000111100001111000010011001100110010110011001100110,
64'b1001011010010110100101101001011010010110011010010110100110010110,
64'b1010010101011010101001010101101001100110100110011001100101100110,
64'b1100110011001100110011001100110000111100001111000011110000111100,
64'b1111111111111111000000000000000011111111000000001111111100000000,
64'b1100110011001100110011001100110001010101101010100101010110101010,
64'b1010010110100101010110100101101001100110100110011001100101100110,
64'b1010010110100101010110100101101010011001100110010110011001100110,
64'b1001100101100110100110010110011000000000000000000000000000000000,
64'b1111111100000000111111110000000000111100110000111100001100111100,
64'b0110011001100110011001100110011010101010101010101010101010101010,
64'b1100110000110011001100111100110010101010010101010101010110101010,
64'b1001100110011001011001100110011010010110100101101001011010010110,
64'b0101010110101010010101011010101000111100001111000011110000111100,
64'b1100001100111100110000110011110010010110011010010110100110010110,
64'b1100110000110011001100111100110001101001011010011001011010010110,
64'b1111000011110000111100001111000010100101010110101010010101011010,
64'b0000000000000000000000000000000011111111111111110000000000000000,
64'b0101101001011010010110100101101000110011001100111100110011001100,
64'b0011001111001100001100111100110011000011110000110011110000111100,
64'b1001100101100110100110010110011010010110100101101001011010010110,
64'b0110100101101001100101101001011010101010101010101010101010101010,
64'b1111111111111111000000000000000011110000000011110000111111110000,
64'b0011110000111100001111000011110001100110011001100110011001100110,
64'b1111000000001111000011111111000000110011001100111100110011001100,
64'b0110100110010110011010011001011001101001100101100110100110010110,
64'b1111000011110000111100001111000000001111111100000000111111110000,
64'b1111111111111111000000000000000000111100110000111100001100111100,
64'b0000000000000000000000000000000001101001100101100110100110010110,
64'b0011001100110011110011001100110001100110100110011001100101100110,
64'b0011110000111100001111000011110000000000000000000000000000000000,
64'b1111000000001111000011111111000001011010010110100101101001011010,
64'b0011110011000011110000110011110010100101010110101010010101011010,
64'b0011001111001100001100111100110001101001100101100110100110010110,
64'b1010010101011010101001010101101011001100110011001100110011001100,
64'b1010101001010101010101011010101000000000111111111111111100000000,
64'b0011110000111100001111000011110010010110100101101001011010010110,
64'b1111111111111111000000000000000001011010010110100101101001011010,
64'b0110100101101001100101101001011010010110011010010110100110010110,
64'b1001011001101001011010011001011000000000111111111111111100000000,
64'b0000111111110000000011111111000011110000000011110000111111110000,
64'b1010010110100101010110100101101010010110011010010110100110010110,
64'b1001011001101001011010011001011011000011110000110011110000111100,
64'b1001100101100110100110010110011010101010101010101010101010101010,
64'b1100001100111100110000110011110000110011110011000011001111001100,
64'b0110100101101001100101101001011011001100001100110011001111001100,
64'b0101010110101010010101011010101000111100110000111100001100111100,
64'b1010101001010101010101011010101011110000111100001111000011110000,
64'b0011001111001100001100111100110011111111111111110000000000000000,
64'b0011110000111100001111000011110001101001100101100110100110010110,
64'b1010101010101010101010101010101001100110011001100110011001100110,
64'b0110100110010110011010011001011011000011110000110011110000111100,
64'b1001011001101001011010011001011000111100001111000011110000111100,
64'b1010101001010101010101011010101010100101101001010101101001011010,
64'b0011001111001100001100111100110010011001011001101001100101100110,
64'b1001011001101001011010011001011011000011110000110011110000111100,
64'b0110100101101001100101101001011001011010010110100101101001011010,
64'b1111000000001111000011111111000011001100110011001100110011001100,
64'b1100001100111100110000110011110000111100110000111100001100111100,
64'b1001100110011001011001100110011010101010101010101010101010101010,
64'b0011001100110011110011001100110000110011110011000011001111001100,
64'b1010010110100101010110100101101000000000111111111111111100000000,
64'b0000111111110000000011111111000011110000111100001111000011110000,
64'b0011001111001100001100111100110001101001100101100110100110010110,
64'b1100001111000011001111000011110011110000111100001111000011110000,
64'b0101010110101010010101011010101011001100001100110011001111001100,
64'b1001011001101001011010011001011000111100001111000011110000111100,
64'b1010101010101010101010101010101001100110011001100110011001100110,
64'b0101101001011010010110100101101001101001011010011001011010010110,
64'b0101010110101010010101011010101010100101010110101010010101011010,
64'b0110100110010110011010011001011000110011001100111100110011001100,
64'b0110100101101001100101101001011011000011110000110011110000111100,
64'b1100110000110011001100111100110010010110011010010110100110010110,
64'b0011110000111100001111000011110001101001011010011001011010010110,
64'b1001100110011001011001100110011011111111000000001111111100000000,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b0101101010100101101001010101101010010110011010010110100110010110,
64'b1111000011110000111100001111000011111111000000001111111100000000,
64'b1111000011110000111100001111000000001111000011111111000011110000,
64'b0011001100110011110011001100110010100101010110101010010101011010,
64'b0110100101101001100101101001011000111100001111000011110000111100,
64'b0101010101010101101010101010101011000011001111001100001100111100,
64'b0000111100001111111100001111000001100110100110011001100101100110,
64'b1111111100000000111111110000000011110000111100001111000011110000,
64'b1111000011110000111100001111000010100101010110101010010101011010,
64'b0101010110101010010101011010101010010110011010010110100110010110,
64'b1100001100111100110000110011110001101001100101100110100110010110,
64'b0011110011000011110000110011110001010101010101011010101010101010,
64'b1100001100111100110000110011110011110000111100001111000011110000,
64'b0110011010011001100110010110011000111100110000111100001100111100,
64'b0101010110101010010101011010101001010101010101011010101010101010,
64'b1111111100000000111111110000000011111111000000001111111100000000,
64'b1111000011110000111100001111000001100110100110011001100101100110,
64'b0110100110010110011010011001011000001111111100000000111111110000,
64'b0110011001100110011001100110011011110000000011110000111111110000,
64'b0101010110101010010101011010101011000011110000110011110000111100,
64'b0101010101010101101010101010101001010101101010100101010110101010,
64'b1111111100000000111111110000000011001100001100110011001111001100,
64'b0011001100110011110011001100110000111100110000111100001100111100,
64'b1111000000001111000011111111000010010110011010010110100110010110,
64'b1111000000001111000011111111000011001100110011001100110011001100,
64'b1010010101011010101001010101101001010101101010100101010110101010,
64'b0011110011000011110000110011110000001111000011111111000011110000,
64'b0110011010011001100110010110011010011001011001101001100101100110,
64'b1001011010010110100101101001011000111100001111000011110000111100,
64'b1111000011110000111100001111000011001100001100110011001111001100,
64'b0011001111001100001100111100110010100101010110101010010101011010,
64'b0101101010100101101001010101101001100110011001100110011001100110,
64'b0000111100001111111100001111000010011001011001101001100101100110,
64'b0000111100001111111100001111000001011010010110100101101001011010,
64'b0110011010011001100110010110011000111100110000111100001100111100,
64'b0000000011111111111111110000000010101010101010101010101010101010,
64'b1100110000110011001100111100110011110000000011110000111111110000,
64'b1010101010101010101010101010101001011010101001011010010101011010,
64'b0000000000000000000000000000000001010101101010100101010110101010,
64'b0000111100001111111100001111000011111111000000001111111100000000,
64'b1001011001101001011010011001011001101001011010011001011010010110,
64'b0000000011111111111111110000000000001111111100000000111111110000,
64'b1111000011110000111100001111000000001111000011111111000011110000,
64'b0000000000000000000000000000000001100110100110011001100101100110,
64'b1010101010101010101010101010101000111100001111000011110000111100,
64'b0110100110010110011010011001011011000011110000110011110000111100,
64'b1001011001101001011010011001011000110011110011000011001111001100,
64'b0101101010100101101001010101101011110000000011110000111111110000,
64'b1010010101011010101001010101101001100110011001100110011001100110,
64'b1100001111000011001111000011110000000000111111111111111100000000,
64'b0110011010011001100110010110011001100110100110011001100101100110,
64'b1001100101100110100110010110011001100110011001100110011001100110,
64'b1010101010101010101010101010101011111111111111110000000000000000,
64'b0110100101101001100101101001011011000011001111001100001100111100,
64'b0011110000111100001111000011110010101010010101010101010110101010,
64'b0101101001011010010110100101101011111111000000001111111100000000,
64'b0000111100001111111100001111000001101001011010011001011010010110,
64'b1010101001010101010101011010101010100101010110101010010101011010,
64'b0000000011111111111111110000000000001111111100000000111111110000,
64'b1111111100000000111111110000000010100101101001010101101001011010,
64'b0101010101010101101010101010101000000000111111111111111100000000,
64'b1001011010010110100101101001011010010110100101101001011010010110,
64'b0110100110010110011010011001011011111111111111110000000000000000,
64'b0110100110010110011010011001011001101001011010011001011010010110,
64'b0000111111110000000011111111000010010110100101101001011010010110,
64'b1100110011001100110011001100110010101010101010101010101010101010,
64'b1100001100111100110000110011110001011010101001011010010101011010,
64'b1010010101011010101001010101101000110011001100111100110011001100,
64'b0011001111001100001100111100110001010101010101011010101010101010,
64'b1111111100000000111111110000000011000011001111001100001100111100,
64'b1001100110011001011001100110011001100110100110011001100101100110,
64'b0101010101010101101010101010101000000000111111111111111100000000,
64'b0101010101010101101010101010101000110011110011000011001111001100,
64'b1100110011001100110011001100110001010101010101011010101010101010,
64'b0110100110010110011010011001011001101001100101100110100110010110,
64'b0011110011000011110000110011110000000000000000000000000000000000,
64'b0011110011000011110000110011110001101001100101100110100110010110,
64'b1111111100000000111111110000000001101001100101100110100110010110,
64'b0101101001011010010110100101101011001100110011001100110011001100,
64'b1111000000001111000011111111000011001100001100110011001111001100,
64'b1100110000110011001100111100110001011010010110100101101001011010,
64'b0000111100001111111100001111000001100110011001100110011001100110,
64'b1111111111111111000000000000000001011010101001011010010101011010,
64'b0011110000111100001111000011110011000011110000110011110000111100,
64'b0110011001100110011001100110011001010101010101011010101010101010,
64'b0110011001100110011001100110011010100101101001010101101001011010,
64'b0101101001011010010110100101101011001100110011001100110011001100,
64'b0011110011000011110000110011110010010110011010010110100110010110,
64'b1111000000001111000011111111000000000000000000000000000000000000,
64'b0101101010100101101001010101101000111100110000111100001100111100,
64'b1010101010101010101010101010101011000011001111001100001100111100,
64'b1001100101100110100110010110011011110000111100001111000011110000,
64'b0000000011111111111111110000000000001111000011111111000011110000,
64'b1010010110100101010110100101101010011001011001101001100101100110,
64'b0101010110101010010101011010101000111100001111000011110000111100,
64'b1010101010101010101010101010101011001100001100110011001111001100,
64'b1010010101011010101001010101101010100101010110101010010101011010,
64'b0011110000111100001111000011110001100110011001100110011001100110,
64'b0011110000111100001111000011110010011001011001101001100101100110,
64'b0011001111001100001100111100110001011010010110100101101001011010,
64'b1111000000001111000011111111000000111100110000111100001100111100,
64'b1010101001010101010101011010101010101010101010101010101010101010,
64'b0110011010011001100110010110011011110000000011110000111111110000,
64'b0110011001100110011001100110011010100101010110101010010101011010,
64'b1001011010010110100101101001011010011001011001101001100101100110,
64'b0101101010100101101001010101101010101010010101010101010110101010,
64'b1001011001101001011010011001011011000011001111001100001100111100,
64'b1001100101100110100110010110011000000000000000000000000000000000,
64'b0101101001011010010110100101101010100101101001010101101001011010,
64'b0101010110101010010101011010101000001111111100000000111111110000,
64'b0101101001011010010110100101101010010110100101101001011010010110,
64'b0101101010100101101001010101101010100101101001010101101001011010,
64'b0000111100001111111100001111000011000011110000110011110000111100,
64'b0000111100001111111100001111000010101010010101010101010110101010,
64'b0101101010100101101001010101101000111100001111000011110000111100,
64'b0000000011111111111111110000000010011001011001101001100101100110,
64'b1010101010101010101010101010101010010110100101101001011010010110,
64'b1111111100000000111111110000000001101001011010011001011010010110,
64'b1001011010010110100101101001011000110011001100111100110011001100,
64'b0000000000000000000000000000000001011010101001011010010101011010,
64'b1111000000001111000011111111000000000000000000000000000000000000,
64'b0110100110010110011010011001011000110011110011000011001111001100,
64'b0110011010011001100110010110011010101010010101010101010110101010,
64'b0110100110010110011010011001011011000011001111001100001100111100,
64'b1001011010010110100101101001011000110011110011000011001111001100,
64'b0101101010100101101001010101101010100101010110101010010101011010,
64'b0101101010100101101001010101101010011001100110010110011001100110,
64'b0011110000111100001111000011110010100101010110101010010101011010,
64'b0101010110101010010101011010101011000011110000110011110000111100,
64'b1100110011001100110011001100110011000011001111001100001100111100,
64'b1100001111000011001111000011110001101001100101100110100110010110,
64'b1001100110011001011001100110011001011010010110100101101001011010,
64'b1001011001101001011010011001011001100110100110011001100101100110,
64'b1001100110011001011001100110011010101010101010101010101010101010,
64'b1100110000110011001100111100110000001111000011111111000011110000,
64'b1001011001101001011010011001011000110011001100111100110011001100,
64'b1100110000110011001100111100110001011010101001011010010101011010,
64'b1001100110011001011001100110011000001111000011111111000011110000,
64'b1100001100111100110000110011110011001100001100110011001111001100,
64'b0110100110010110011010011001011000111100001111000011110000111100,
64'b1111111111111111000000000000000001100110100110011001100101100110,
64'b0011001111001100001100111100110000001111111100000000111111110000,
64'b0101101001011010010110100101101010100101010110101010010101011010,
64'b0000111111110000000011111111000000111100110000111100001100111100,
64'b1001011010010110100101101001011000110011110011000011001111001100,
64'b1001011001101001011010011001011011000011110000110011110000111100,
64'b1001011010010110100101101001011001100110011001100110011001100110,
64'b1010010110100101010110100101101011111111000000001111111100000000,
64'b1001011001101001011010011001011001011010010110100101101001011010,
64'b1010010110100101010110100101101001100110100110011001100101100110,
64'b1001011010010110100101101001011001010101101010100101010110101010,
64'b0101101010100101101001010101101010100101101001010101101001011010,
64'b0011110011000011110000110011110010100101010110101010010101011010,
64'b0000000000000000000000000000000011000011110000110011110000111100,
64'b1010010110100101010110100101101010101010010101010101010110101010,
64'b0011001111001100001100111100110000110011110011000011001111001100,
64'b1001011001101001011010011001011011110000000011110000111111110000,
64'b1001100110011001011001100110011010100101101001010101101001011010,
64'b1010101010101010101010101010101000001111111100000000111111110000,
64'b1111000011110000111100001111000010010110100101101001011010010110,
64'b0110100110010110011010011001011011111111111111110000000000000000,
64'b1100001111000011001111000011110000110011110011000011001111001100,
64'b1100001100111100110000110011110011000011110000110011110000111100,
64'b0011001100110011110011001100110010011001100110010110011001100110,
64'b1100001100111100110000110011110000110011110011000011001111001100,
64'b0101010110101010010101011010101001100110100110011001100101100110,
64'b1111000000001111000011111111000000001111111100000000111111110000,
64'b0011001100110011110011001100110010011001100110010110011001100110,
64'b1111000011110000111100001111000001011010010110100101101001011010,
64'b1010101001010101010101011010101000000000111111111111111100000000,
64'b1100110000110011001100111100110010011001011001101001100101100110,
64'b1111000000001111000011111111000010101010010101010101010110101010,
64'b0110011001100110011001100110011011000011001111001100001100111100,
64'b0110011010011001100110010110011000000000000000000000000000000000,
64'b0101101001011010010110100101101010100101101001010101101001011010,
64'b0000000011111111111111110000000000001111111100000000111111110000,
64'b1010101001010101010101011010101010010110100101101001011010010110,
64'b0101010110101010010101011010101010100101101001010101101001011010,
64'b0011110000111100001111000011110011000011110000110011110000111100,
64'b0101101001011010010110100101101010101010010101010101010110101010,
64'b0101101010100101101001010101101000111100001111000011110000111100,
64'b1111111100000000111111110000000010011001011001101001100101100110,
64'b0011001100110011110011001100110011000011110000110011110000111100,
64'b1010010110100101010110100101101000110011110011000011001111001100,
64'b1010101001010101010101011010101010100101010110101010010101011010,
64'b1001011010010110100101101001011011000011110000110011110000111100,
64'b1100001111000011001111000011110001011010010110100101101001011010,
64'b1001100101100110100110010110011001100110011001100110011001100110,
64'b1111111111111111000000000000000011110000000011110000111111110000,
64'b1001100110011001011001100110011010011001100110010110011001100110,
64'b1001100110011001011001100110011000111100110000111100001100111100,
64'b0000111111110000000011111111000010101010010101010101010110101010,
64'b0011001111001100001100111100110011000011001111001100001100111100,
64'b1100110000110011001100111100110010100101101001010101101001011010,
64'b1010101010101010101010101010101010010110100101101001011010010110,
64'b1100110011001100110011001100110010011001011001101001100101100110,
64'b1100001111000011001111000011110011111111000000001111111100000000,
64'b0000111111110000000011111111000001011010010110100101101001011010,
64'b1111000011110000111100001111000010010110100101101001011010010110,
64'b0101010110101010010101011010101011000011001111001100001100111100,
64'b0011110011000011110000110011110001101001100101100110100110010110,
64'b0101101001011010010110100101101001011010101001011010010101011010,
64'b1100110000110011001100111100110011001100001100110011001111001100,
64'b1001100110011001011001100110011001010101101010100101010110101010,
64'b1010010101011010101001010101101010010110100101101001011010010110,
64'b0101010110101010010101011010101000000000000000000000000000000000,
64'b0000111111110000000011111111000000110011001100111100110011001100,
64'b1100110011001100110011001100110011000011001111001100001100111100,
64'b0110011001100110011001100110011011000011110000110011110000111100,
64'b0101010101010101101010101010101011111111111111110000000000000000,
64'b0011110000111100001111000011110000110011110011000011001111001100,
64'b0110011001100110011001100110011011000011001111001100001100111100,
64'b0110100101101001100101101001011011110000000011110000111111110000,
64'b1010010110100101010110100101101000111100110000111100001100111100,
64'b1100001100111100110000110011110011001100001100110011001111001100,
64'b0101010110101010010101011010101010100101101001010101101001011010,
64'b1001100110011001011001100110011010011001100110010110011001100110,
64'b0110100110010110011010011001011011000011001111001100001100111100,
64'b0110100110010110011010011001011000000000000000000000000000000000,
64'b0000000000000000000000000000000011110000111100001111000011110000,
64'b0101101001011010010110100101101010100101010110101010010101011010,
64'b1001011010010110100101101001011000001111111100000000111111110000,
64'b1100110011001100110011001100110010101010101010101010101010101010,
64'b1010010101011010101001010101101010100101101001010101101001011010,
64'b0011110000111100001111000011110011110000000011110000111111110000,
64'b1100001100111100110000110011110000000000111111111111111100000000,
64'b1001100101100110100110010110011001011010101001011010010101011010,
64'b0101101010100101101001010101101010100101101001010101101001011010,
64'b0011001100110011110011001100110010011001011001101001100101100110,
64'b0011110000111100001111000011110010010110100101101001011010010110,
64'b1001011001101001011010011001011001011010101001011010010101011010,
64'b0011110011000011110000110011110000000000000000000000000000000000,
64'b0000000000000000000000000000000011111111000000001111111100000000,
64'b0011001111001100001100111100110000110011110011000011001111001100,
64'b1111111100000000111111110000000000111100110000111100001100111100,
64'b1010101001010101010101011010101010010110011010010110100110010110,
64'b0101101001011010010110100101101010100101101001010101101001011010,
64'b1001011010010110100101101001011000110011001100111100110011001100,
64'b1010101001010101010101011010101000001111000011111111000011110000,
64'b1001011001101001011010011001011000110011001100111100110011001100,
64'b1001011001101001011010011001011011000011001111001100001100111100,
64'b0000000011111111111111110000000000110011110011000011001111001100,
64'b1010101001010101010101011010101011001100001100110011001111001100,
64'b0011001111001100001100111100110011000011001111001100001100111100,
64'b0000000000000000000000000000000011110000000011110000111111110000,
64'b1010101001010101010101011010101011111111000000001111111100000000,
64'b0101101001011010010110100101101001011010010110100101101001011010,
64'b0110100101101001100101101001011001011010101001011010010101011010,
64'b0110100110010110011010011001011010010110011010010110100110010110,
64'b0000111100001111111100001111000010011001011001101001100101100110,
64'b0101101001011010010110100101101001011010010110100101101001011010,
64'b0110100101101001100101101001011001010101101010100101010110101010,
64'b1100001111000011001111000011110001011010010110100101101001011010,
64'b1100110000110011001100111100110001011010101001011010010101011010,
64'b0000111111110000000011111111000000001111000011111111000011110000,
64'b1001011010010110100101101001011000001111000011111111000011110000,
64'b1010101010101010101010101010101001011010101001011010010101011010,
64'b0101101010100101101001010101101000000000111111111111111100000000,
64'b0011001111001100001100111100110001010101010101011010101010101010,
64'b0011001111001100001100111100110000110011110011000011001111001100,
64'b1111111100000000111111110000000011001100001100110011001111001100,
64'b1100110011001100110011001100110010010110011010010110100110010110,
64'b0110100101101001100101101001011001101001011010011001011010010110,
64'b0000000000000000000000000000000000110011110011000011001111001100,
64'b1001100101100110100110010110011000110011001100111100110011001100,
64'b1111000011110000111100001111000000110011110011000011001111001100,
64'b1111111111111111000000000000000011001100001100110011001111001100,
64'b1111000011110000111100001111000001010101101010100101010110101010,
64'b1100110000110011001100111100110001010101101010100101010110101010,
64'b1100001111000011001111000011110001100110100110011001100101100110,
64'b1001011010010110100101101001011001010101010101011010101010101010,
64'b1010010101011010101001010101101001100110011001100110011001100110,
64'b0101101001011010010110100101101001011010010110100101101001011010,
64'b0101010101010101101010101010101000001111000011111111000011110000,
64'b1111000011110000111100001111000010010110011010010110100110010110,
64'b1100001100111100110000110011110001101001100101100110100110010110,
64'b1010101010101010101010101010101010100101101001010101101001011010,
64'b1100001111000011001111000011110011110000111100001111000011110000,
64'b1111111100000000111111110000000010100101101001010101101001011010,
64'b0000000000000000000000000000000000001111000011111111000011110000,
64'b0101010110101010010101011010101010011001100110010110011001100110,
64'b0000111100001111111100001111000000110011001100111100110011001100,
64'b1010010101011010101001010101101011000011110000110011110000111100,
64'b0110100110010110011010011001011001100110011001100110011001100110,
64'b1100110000110011001100111100110010010110100101101001011010010110,
64'b0011001111001100001100111100110000110011110011000011001111001100,
64'b0110011001100110011001100110011001010101101010100101010110101010,
64'b0101010110101010010101011010101010010110011010010110100110010110,
64'b1111000000001111000011111111000010010110011010010110100110010110,
64'b1100110011001100110011001100110000110011110011000011001111001100,
64'b0000111111110000000011111111000001010101101010100101010110101010,
64'b0101010101010101101010101010101000110011110011000011001111001100,
64'b0000000000000000000000000000000001010101101010100101010110101010,
64'b0011001100110011110011001100110010010110100101101001011010010110,
64'b1111111100000000111111110000000001011010010110100101101001011010,
64'b0110011010011001100110010110011010100101010110101010010101011010,
64'b0011110011000011110000110011110010010110100101101001011010010110,
64'b0000111100001111111100001111000011000011001111001100001100111100,
64'b0101101001011010010110100101101011110000111100001111000011110000,
64'b0011110000111100001111000011110010011001100110010110011001100110,
64'b0011001100110011110011001100110000111100110000111100001100111100,
64'b0000000011111111111111110000000010010110011010010110100110010110,
64'b0101101001011010010110100101101010100101101001010101101001011010,
64'b0000000011111111111111110000000000110011001100111100110011001100,
64'b1100110011001100110011001100110000001111000011111111000011110000,
64'b1010101010101010101010101010101000110011001100111100110011001100,
64'b1111000011110000111100001111000011000011001111001100001100111100,
64'b0101010101010101101010101010101000110011110011000011001111001100,
64'b1100001111000011001111000011110011001100001100110011001111001100,
64'b0101101010100101101001010101101011000011001111001100001100111100,
64'b0101010110101010010101011010101011110000000011110000111111110000,
64'b1001100101100110100110010110011011111111000000001111111100000000,
64'b1010010110100101010110100101101011111111111111110000000000000000,
64'b0000111100001111111100001111000001100110100110011001100101100110,
64'b1001100101100110100110010110011011111111000000001111111100000000,
64'b1010101001010101010101011010101010101010010101010101010110101010,
64'b0110011010011001100110010110011010100101010110101010010101011010,
64'b0110011001100110011001100110011011000011001111001100001100111100,
64'b1001100110011001011001100110011000110011110011000011001111001100,
64'b0110100110010110011010011001011010011001100110010110011001100110,
64'b0101010110101010010101011010101000001111000011111111000011110000,
64'b0011110011000011110000110011110011111111111111110000000000000000,
64'b0110100101101001100101101001011000001111111100000000111111110000,
64'b1001011010010110100101101001011000111100110000111100001100111100,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b1001011001101001011010011001011000000000000000000000000000000000,
64'b0101101010100101101001010101101001101001011010011001011010010110,
64'b1111000000001111000011111111000001010101010101011010101010101010,
64'b1001100101100110100110010110011000110011001100111100110011001100,
64'b0000111111110000000011111111000001100110100110011001100101100110,
64'b1111000011110000111100001111000011110000000011110000111111110000,
64'b1010010110100101010110100101101000001111000011111111000011110000,
64'b1111111111111111000000000000000000111100001111000011110000111100,
64'b0110011010011001100110010110011001010101101010100101010110101010,
64'b1100110011001100110011001100110010101010101010101010101010101010,
64'b0000000011111111111111110000000010101010010101010101010110101010,
64'b1111111100000000111111110000000011110000000011110000111111110000,
64'b0011110000111100001111000011110001011010010110100101101001011010,
64'b1001100101100110100110010110011010101010101010101010101010101010,
64'b0110100110010110011010011001011011000011001111001100001100111100,
64'b0011001100110011110011001100110001100110011001100110011001100110,
64'b1100001100111100110000110011110001011010010110100101101001011010,
64'b0110011001100110011001100110011001101001011010011001011010010110,
64'b1001100101100110100110010110011010101010010101010101010110101010,
64'b1010101001010101010101011010101001010101101010100101010110101010,
64'b1100001100111100110000110011110010100101010110101010010101011010,
64'b0011110011000011110000110011110000110011001100111100110011001100,
64'b0110011010011001100110010110011011001100110011001100110011001100,
64'b1001011010010110100101101001011000110011001100111100110011001100,
64'b1100001111000011001111000011110010101010010101010101010110101010,
64'b1100001100111100110000110011110010011001011001101001100101100110,
64'b1100001111000011001111000011110001100110011001100110011001100110,
64'b0011110011000011110000110011110011110000000011110000111111110000,
64'b1111000011110000111100001111000000111100001111000011110000111100,
64'b0101101010100101101001010101101000110011110011000011001111001100,
64'b0011110000111100001111000011110011000011001111001100001100111100,
64'b1100001111000011001111000011110010011001100110010110011001100110,
64'b0011001100110011110011001100110010011001100110010110011001100110,
64'b0101101010100101101001010101101011001100001100110011001111001100,
64'b1111000000001111000011111111000011110000111100001111000011110000,
64'b0110100101101001100101101001011001011010010110100101101001011010,
64'b0110100110010110011010011001011011110000111100001111000011110000,
64'b0000111111110000000011111111000010011001100110010110011001100110,
64'b1010010101011010101001010101101010010110100101101001011010010110,
64'b0000000011111111111111110000000010010110100101101001011010010110,
64'b0101010110101010010101011010101000000000111111111111111100000000,
64'b1100110011001100110011001100110010100101010110101010010101011010,
64'b0110011001100110011001100110011000001111000011111111000011110000,
64'b1100001111000011001111000011110011110000000011110000111111110000,
64'b0110100110010110011010011001011000111100001111000011110000111100,
64'b1100001111000011001111000011110010010110100101101001011010010110,
64'b0000111100001111111100001111000010100101101001010101101001011010,
64'b1111111111111111000000000000000001010101101010100101010110101010,
64'b0101010101010101101010101010101000110011110011000011001111001100,
64'b1111111100000000111111110000000011111111000000001111111100000000,
64'b1001011001101001011010011001011000111100001111000011110000111100,
64'b1111111100000000111111110000000001101001100101100110100110010110,
64'b0101101001011010010110100101101011000011001111001100001100111100,
64'b1001011010010110100101101001011011111111111111110000000000000000,
64'b0110100110010110011010011001011001100110100110011001100101100110,
64'b1001011001101001011010011001011011111111000000001111111100000000,
64'b0110100101101001100101101001011010101010010101010101010110101010,
64'b1111000000001111000011111111000010100101010110101010010101011010,
64'b1001011001101001011010011001011011000011001111001100001100111100,
64'b0011110000111100001111000011110000110011110011000011001111001100,
64'b1111111100000000111111110000000010011001100110010110011001100110,
64'b0101101010100101101001010101101000001111000011111111000011110000,
64'b0011110000111100001111000011110011111111111111110000000000000000,
64'b1010101001010101010101011010101000001111111100000000111111110000,
64'b0110011001100110011001100110011011000011001111001100001100111100,
64'b1001100101100110100110010110011011111111000000001111111100000000,
64'b1100001100111100110000110011110000001111000011111111000011110000,
64'b0011110011000011110000110011110011110000000011110000111111110000,
64'b0011110011000011110000110011110011111111000000001111111100000000,
64'b0110100110010110011010011001011001010101101010100101010110101010,
64'b1010101001010101010101011010101000000000111111111111111100000000,
64'b1001011001101001011010011001011001101001100101100110100110010110,
64'b1010010101011010101001010101101001100110100110011001100101100110,
64'b1111111111111111000000000000000001101001100101100110100110010110,
64'b1100110000110011001100111100110001101001011010011001011010010110,
64'b1010010101011010101001010101101011000011110000110011110000111100,
64'b0011001100110011110011001100110000111100110000111100001100111100,
64'b1001011010010110100101101001011011000011001111001100001100111100,
64'b0110011001100110011001100110011001011010010110100101101001011010,
64'b1111111100000000111111110000000011110000000011110000111111110000,
64'b0110100101101001100101101001011000110011001100111100110011001100,
64'b1111000011110000111100001111000011111111000000001111111100000000,
64'b1111000011110000111100001111000001010101101010100101010110101010,
64'b0101010101010101101010101010101010011001100110010110011001100110,
64'b0000111111110000000011111111000000001111111100000000111111110000,
64'b0000111100001111111100001111000010101010010101010101010110101010,
64'b0101010110101010010101011010101011000011110000110011110000111100,
64'b1001100101100110100110010110011011111111111111110000000000000000,
64'b0000111111110000000011111111000011001100001100110011001111001100,
64'b0110011001100110011001100110011011001100001100110011001111001100,
64'b1010010101011010101001010101101001101001100101100110100110010110,
64'b1001100110011001011001100110011010011001011001101001100101100110,
64'b1111000011110000111100001111000000000000111111111111111100000000,
64'b0101101001011010010110100101101001011010010110100101101001011010,
64'b1111111111111111000000000000000001010101010101011010101010101010,
64'b1001100110011001011001100110011000110011001100111100110011001100,
64'b1010101010101010101010101010101000111100001111000011110000111100,
64'b0011001111001100001100111100110010101010010101010101010110101010,
64'b1001011010010110100101101001011000110011001100111100110011001100,
64'b1100110000110011001100111100110010100101010110101010010101011010,
64'b1111111100000000111111110000000010101010101010101010101010101010,
64'b0110100110010110011010011001011010100101101001010101101001011010,
64'b1010101010101010101010101010101010100101101001010101101001011010,
64'b1111111100000000111111110000000001101001100101100110100110010110,
64'b0011110000111100001111000011110001101001011010011001011010010110,
64'b0101010110101010010101011010101011111111111111110000000000000000,
64'b0011001111001100001100111100110010011001011001101001100101100110,
64'b0000000000000000000000000000000011001100110011001100110011001100,
64'b1001011010010110100101101001011001011010010110100101101001011010,
64'b0110011001100110011001100110011010100101010110101010010101011010,
64'b0000111100001111111100001111000000110011001100111100110011001100,
64'b1100001100111100110000110011110001011010010110100101101001011010,
64'b0000111100001111111100001111000001100110100110011001100101100110,
64'b0101010101010101101010101010101011001100110011001100110011001100,
64'b0011110011000011110000110011110000110011110011000011001111001100,
64'b1100110011001100110011001100110010011001011001101001100101100110,
64'b0000000000000000000000000000000001101001100101100110100110010110,
64'b0000000011111111111111110000000011001100001100110011001111001100,
64'b0011110000111100001111000011110010100101101001010101101001011010,
64'b1001011001101001011010011001011011110000000011110000111111110000,
64'b1010101001010101010101011010101001011010101001011010010101011010,
64'b1010010110100101010110100101101001010101010101011010101010101010,
64'b0101101001011010010110100101101010101010010101010101010110101010,
64'b0110011010011001100110010110011001101001011010011001011010010110,
64'b0011001100110011110011001100110011110000111100001111000011110000,
64'b1010101010101010101010101010101010010110011010010110100110010110,
64'b0101101010100101101001010101101001100110100110011001100101100110,
64'b0011001111001100001100111100110001100110011001100110011001100110,
64'b1100110011001100110011001100110001010101010101011010101010101010,
64'b1100110011001100110011001100110000001111111100000000111111110000,
64'b0101101001011010010110100101101000001111000011111111000011110000,
64'b1010101001010101010101011010101010011001011001101001100101100110,
64'b1010010110100101010110100101101010101010010101010101010110101010,
64'b0011001111001100001100111100110001100110100110011001100101100110,
64'b1111111111111111000000000000000001100110011001100110011001100110,
64'b1111111100000000111111110000000010011001100110010110011001100110,
64'b0101101001011010010110100101101001101001100101100110100110010110,
64'b0011001111001100001100111100110001010101101010100101010110101010,
64'b0011001111001100001100111100110000111100110000111100001100111100,
64'b1111000011110000111100001111000001101001011010011001011010010110,
64'b1100110011001100110011001100110010010110100101101001011010010110,
64'b0110011001100110011001100110011011001100110011001100110011001100,
64'b0011110000111100001111000011110001010101101010100101010110101010,
64'b0011110011000011110000110011110001010101101010100101010110101010,
64'b0011110000111100001111000011110001101001011010011001011010010110,
64'b0000000000000000000000000000000000110011001100111100110011001100,
64'b0000111111110000000011111111000001101001011010011001011010010110,
64'b0110011010011001100110010110011010010110100101101001011010010110,
64'b0011001100110011110011001100110000111100001111000011110000111100,
64'b1010101001010101010101011010101010010110011010010110100110010110,
64'b0110011010011001100110010110011000110011001100111100110011001100,
64'b0101101010100101101001010101101011110000000011110000111111110000,
64'b1100001111000011001111000011110001101001100101100110100110010110,
64'b1001100110011001011001100110011001101001100101100110100110010110,
64'b1010101010101010101010101010101011110000111100001111000011110000,
64'b1100001100111100110000110011110011001100110011001100110011001100,
64'b1111000000001111000011111111000000110011001100111100110011001100,
64'b1010010101011010101001010101101011000011001111001100001100111100,
64'b0000000000000000000000000000000001011010010110100101101001011010,
64'b0000000011111111111111110000000001101001100101100110100110010110,
64'b1100001111000011001111000011110001101001100101100110100110010110,
64'b0101101001011010010110100101101000001111111100000000111111110000,
64'b1001100110011001011001100110011000111100110000111100001100111100,
64'b0110100101101001100101101001011001011010010110100101101001011010,
64'b0110011010011001100110010110011010101010010101010101010110101010,
64'b1010010101011010101001010101101010010110011010010110100110010110,
64'b1001011010010110100101101001011000111100110000111100001100111100,
64'b0110011001100110011001100110011011111111000000001111111100000000,
64'b0000111111110000000011111111000011110000111100001111000011110000,
64'b1010101001010101010101011010101001011010010110100101101001011010,
64'b0110011010011001100110010110011001011010101001011010010101011010,
64'b0000000000000000000000000000000000110011110011000011001111001100,
64'b1111111111111111000000000000000000111100110000111100001100111100,
64'b1010010101011010101001010101101000111100110000111100001100111100,
64'b1001100101100110100110010110011000000000111111111111111100000000,
64'b0011110000111100001111000011110011110000000011110000111111110000,
64'b0110100110010110011010011001011010011001011001101001100101100110,
64'b0110100101101001100101101001011000110011001100111100110011001100,
64'b0110011010011001100110010110011010010110011010010110100110010110,
64'b1100001100111100110000110011110001011010101001011010010101011010,
64'b0011110000111100001111000011110001010101010101011010101010101010,
64'b1111111100000000111111110000000011111111000000001111111100000000,
64'b0011001100110011110011001100110000110011110011000011001111001100,
64'b0110100101101001100101101001011011001100001100110011001111001100,
64'b1010101010101010101010101010101010100101101001010101101001011010,
64'b0000000000000000000000000000000011110000000011110000111111110000,
64'b0110011010011001100110010110011001011010101001011010010101011010,
64'b1100001111000011001111000011110001010101010101011010101010101010,
64'b0000111111110000000011111111000010101010010101010101010110101010,
64'b0011110011000011110000110011110001101001011010011001011010010110,
64'b1100001100111100110000110011110011110000111100001111000011110000,
64'b0110100101101001100101101001011010010110011010010110100110010110,
64'b0101101010100101101001010101101001100110100110011001100101100110,
64'b0000111111110000000011111111000001100110011001100110011001100110,
64'b0000000000000000000000000000000010101010101010101010101010101010,
64'b0011001100110011110011001100110011110000000011110000111111110000,
64'b0110011010011001100110010110011011111111000000001111111100000000,
64'b0110100101101001100101101001011010101010101010101010101010101010,
64'b0101010101010101101010101010101010010110100101101001011010010110,
64'b0011110011000011110000110011110010011001100110010110011001100110,
64'b0011110000111100001111000011110011111111111111110000000000000000,
64'b0011001100110011110011001100110010010110011010010110100110010110,
64'b1001011010010110100101101001011000000000000000000000000000000000,
64'b0101101001011010010110100101101010010110011010010110100110010110,
64'b1010101010101010101010101010101000000000111111111111111100000000,
64'b0000111100001111111100001111000001010101101010100101010110101010,
64'b0110100101101001100101101001011000110011110011000011001111001100,
64'b0000000000000000000000000000000001101001100101100110100110010110,
64'b1100001111000011001111000011110000000000111111111111111100000000,
64'b0000111111110000000011111111000001010101010101011010101010101010,
64'b0000000011111111111111110000000011001100110011001100110011001100,
64'b0011001100110011110011001100110011000011001111001100001100111100,
64'b0110011001100110011001100110011000111100001111000011110000111100,
64'b1001100101100110100110010110011010101010101010101010101010101010,
64'b1100001111000011001111000011110010010110011010010110100110010110,
64'b1111111100000000111111110000000010101010101010101010101010101010,
64'b0110100110010110011010011001011000111100110000111100001100111100,
64'b0110011001100110011001100110011001010101010101011010101010101010,
64'b1111000000001111000011111111000010011001100110010110011001100110,
64'b0000000011111111111111110000000000001111000011111111000011110000,
64'b1010101010101010101010101010101011000011001111001100001100111100,
64'b0011110011000011110000110011110011111111111111110000000000000000,
64'b1100110011001100110011001100110001100110011001100110011001100110,
64'b1001011010010110100101101001011001011010010110100101101001011010,
64'b0000111100001111111100001111000011110000000011110000111111110000,
64'b1010101001010101010101011010101000001111111100000000111111110000,
64'b1111111111111111000000000000000011001100110011001100110011001100,
64'b0011110011000011110000110011110000111100110000111100001100111100,
64'b1100001111000011001111000011110001100110011001100110011001100110,
64'b0110011010011001100110010110011011110000000011110000111111110000,
64'b1001011010010110100101101001011001100110011001100110011001100110,
64'b0000111111110000000011111111000010010110100101101001011010010110,
64'b0011110000111100001111000011110001010101101010100101010110101010,
64'b0110011001100110011001100110011010100101010110101010010101011010,
64'b0101101010100101101001010101101010101010101010101010101010101010,
64'b0101101001011010010110100101101010010110100101101001011010010110,
64'b1100001100111100110000110011110000110011110011000011001111001100,
64'b1111111100000000111111110000000000000000111111111111111100000000,
64'b1001100110011001011001100110011010101010010101010101010110101010,
64'b1010101010101010101010101010101011110000111100001111000011110000,
64'b0101101010100101101001010101101011110000000011110000111111110000,
64'b1010010101011010101001010101101010010110100101101001011010010110,
64'b0110100101101001100101101001011000000000111111111111111100000000,
64'b0110100110010110011010011001011010010110100101101001011010010110,
64'b0000000011111111111111110000000011000011001111001100001100111100,
64'b0000111111110000000011111111000000110011001100111100110011001100,
64'b0011110000111100001111000011110000110011110011000011001111001100,
64'b0101010110101010010101011010101011001100110011001100110011001100,
64'b1111111111111111000000000000000011000011001111001100001100111100,
64'b1001100101100110100110010110011000001111000011111111000011110000,
64'b1010101010101010101010101010101011111111111111110000000000000000,
64'b0000000011111111111111110000000010011001100110010110011001100110,
64'b0101101001011010010110100101101001010101101010100101010110101010,
64'b1111111100000000111111110000000000000000111111111111111100000000,
64'b1111000000001111000011111111000001101001100101100110100110010110,
64'b1001100101100110100110010110011011111111111111110000000000000000,
64'b0011110011000011110000110011110001101001100101100110100110010110,
64'b1111000011110000111100001111000011110000000011110000111111110000,
64'b1100001100111100110000110011110011110000111100001111000011110000,
64'b0000111111110000000011111111000001011010010110100101101001011010,
64'b1010101010101010101010101010101001011010010110100101101001011010,
64'b0110011010011001100110010110011011110000000011110000111111110000,
64'b0000000000000000000000000000000011111111000000001111111100000000,
64'b1001100110011001011001100110011010101010101010101010101010101010,
64'b1100001100111100110000110011110010010110100101101001011010010110,
64'b1010010101011010101001010101101010011001100110010110011001100110,
64'b1100110011001100110011001100110011111111111111110000000000000000,
64'b1001011001101001011010011001011010010110011010010110100110010110,
64'b0011001100110011110011001100110000000000000000000000000000000000,
64'b0101101010100101101001010101101010010110011010010110100110010110,
64'b0101101010100101101001010101101000000000111111111111111100000000,
64'b1001100101100110100110010110011001010101101010100101010110101010,
64'b1111111100000000111111110000000000110011110011000011001111001100,
64'b1100110011001100110011001100110010101010010101010101010110101010,
64'b1100001111000011001111000011110001100110011001100110011001100110,
64'b1010101010101010101010101010101000111100001111000011110000111100,
64'b0011110000111100001111000011110010011001100110010110011001100110,
64'b0101101010100101101001010101101011111111111111110000000000000000,
64'b1100110000110011001100111100110000000000000000000000000000000000,
64'b1111000011110000111100001111000010011001100110010110011001100110,
64'b0011110011000011110000110011110000000000111111111111111100000000,
64'b0101101001011010010110100101101011110000111100001111000011110000,
64'b0110011010011001100110010110011010010110011010010110100110010110,
64'b0110011010011001100110010110011001011010010110100101101001011010,
64'b0110100101101001100101101001011011110000111100001111000011110000,
64'b0000000000000000000000000000000011110000111100001111000011110000,
64'b1100001111000011001111000011110010101010101010101010101010101010,
64'b0110100101101001100101101001011011110000000011110000111111110000,
64'b0000111100001111111100001111000001100110100110011001100101100110,
64'b0101101010100101101001010101101001101001011010011001011010010110,
64'b1111000011110000111100001111000010010110011010010110100110010110,
64'b1001100110011001011001100110011010010110100101101001011010010110,
64'b0110011010011001100110010110011000001111000011111111000011110000,
64'b0110011010011001100110010110011011000011110000110011110000111100,
64'b1100001100111100110000110011110000001111111100000000111111110000,
64'b0110100101101001100101101001011010010110011010010110100110010110,
64'b0110011001100110011001100110011010010110011010010110100110010110,
64'b0000000011111111111111110000000010010110011010010110100110010110,
64'b1010101010101010101010101010101011111111000000001111111100000000,
64'b1001011001101001011010011001011001100110011001100110011001100110,
64'b0000111100001111111100001111000000000000111111111111111100000000,
64'b0011110011000011110000110011110001101001011010011001011010010110,
64'b0011001111001100001100111100110001101001100101100110100110010110,
64'b0110100101101001100101101001011010010110011010010110100110010110,
64'b0000000000000000000000000000000001101001100101100110100110010110,
64'b0101101001011010010110100101101011111111000000001111111100000000,
64'b1111111111111111000000000000000010100101010110101010010101011010,
64'b0000000011111111111111110000000010101010010101010101010110101010,
64'b0110100110010110011010011001011000111100110000111100001100111100,
64'b1001100110011001011001100110011010010110011010010110100110010110,
64'b1001011010010110100101101001011010010110011010010110100110010110,
64'b0110011001100110011001100110011010101010101010101010101010101010,
64'b1001011001101001011010011001011010010110100101101001011010010110,
64'b0101010110101010010101011010101011111111111111110000000000000000,
64'b0101101010100101101001010101101001101001100101100110100110010110,
64'b1010010110100101010110100101101010010110011010010110100110010110,
64'b1100001100111100110000110011110000111100110000111100001100111100,
64'b1010101010101010101010101010101010010110011010010110100110010110,
64'b0011001111001100001100111100110011111111111111110000000000000000,
64'b0000000000000000000000000000000011001100001100110011001111001100,
64'b0101010101010101101010101010101000110011001100111100110011001100,
64'b1001011001101001011010011001011001011010101001011010010101011010,
64'b0011110000111100001111000011110010010110011010010110100110010110,
64'b0110100110010110011010011001011010010110011010010110100110010110,
64'b0011110000111100001111000011110001100110011001100110011001100110,
64'b0000111111110000000011111111000001011010101001011010010101011010,
64'b1111111100000000111111110000000001100110100110011001100101100110,
64'b1010010101011010101001010101101011111111000000001111111100000000,
64'b1100110000110011001100111100110001101001100101100110100110010110,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b1111000011110000111100001111000010101010010101010101010110101010,
64'b0011110000111100001111000011110010011001100110010110011001100110,
64'b1001011010010110100101101001011000110011001100111100110011001100,
64'b1001011010010110100101101001011000000000000000000000000000000000,
64'b0011110011000011110000110011110011001100001100110011001111001100,
64'b1010101001010101010101011010101010011001011001101001100101100110,
64'b0101010110101010010101011010101011111111000000001111111100000000,
64'b0000111111110000000011111111000010010110100101101001011010010110,
64'b0011001111001100001100111100110001100110100110011001100101100110,
64'b1001100101100110100110010110011001101001011010011001011010010110,
64'b1010010101011010101001010101101001010101010101011010101010101010,
64'b0101101001011010010110100101101000111100110000111100001100111100,
64'b1010101001010101010101011010101000111100001111000011110000111100,
64'b1100001100111100110000110011110000110011001100111100110011001100,
64'b0011110011000011110000110011110010010110100101101001011010010110,
64'b0101010110101010010101011010101001011010010110100101101001011010,
64'b1001100101100110100110010110011010101010101010101010101010101010,
64'b0101101010100101101001010101101000001111000011111111000011110000,
64'b1001011010010110100101101001011001101001011010011001011010010110,
64'b1111000011110000111100001111000011111111111111110000000000000000,
64'b1111111100000000111111110000000011000011001111001100001100111100,
64'b0011110000111100001111000011110001101001011010011001011010010110,
64'b1010010101011010101001010101101001101001100101100110100110010110,
64'b1010010101011010101001010101101001100110011001100110011001100110,
64'b0110011010011001100110010110011001011010101001011010010101011010,
64'b0000111111110000000011111111000010100101010110101010010101011010,
64'b0110011010011001100110010110011011110000111100001111000011110000,
64'b1100001100111100110000110011110001101001100101100110100110010110,
64'b0000111100001111111100001111000000110011110011000011001111001100,
64'b1001100110011001011001100110011011001100110011001100110011001100,
64'b0110011010011001100110010110011011111111000000001111111100000000,
64'b0110011010011001100110010110011001101001100101100110100110010110,
64'b1001011001101001011010011001011010101010101010101010101010101010,
64'b0000000000000000000000000000000010100101010110101010010101011010,
64'b1010010101011010101001010101101011000011001111001100001100111100,
64'b1100110000110011001100111100110010010110011010010110100110010110,
64'b1100110000110011001100111100110000111100001111000011110000111100,
64'b1100001111000011001111000011110011001100001100110011001111001100,
64'b1010101001010101010101011010101001100110100110011001100101100110,
64'b1100001111000011001111000011110011111111000000001111111100000000,
64'b0101101010100101101001010101101000111100110000111100001100111100,
64'b1111111100000000111111110000000000001111000011111111000011110000,
64'b1001011010010110100101101001011011110000111100001111000011110000,
64'b0110100101101001100101101001011011111111111111110000000000000000,
64'b0110100101101001100101101001011000111100110000111100001100111100,
64'b1001011001101001011010011001011011001100110011001100110011001100,
64'b1010101010101010101010101010101000110011110011000011001111001100,
64'b0110011010011001100110010110011011110000000011110000111111110000,
64'b0000111100001111111100001111000000111100110000111100001100111100,
64'b1010010110100101010110100101101010100101010110101010010101011010,
64'b1010010101011010101001010101101000001111000011111111000011110000,
64'b1001100110011001011001100110011001101001011010011001011010010110,
64'b1010010101011010101001010101101001010101010101011010101010101010,
64'b0110011010011001100110010110011011110000000011110000111111110000,
64'b0101010101010101101010101010101001010101101010100101010110101010,
64'b1100001100111100110000110011110001010101101010100101010110101010,
64'b1100001100111100110000110011110000000000000000000000000000000000,
64'b0110100110010110011010011001011001011010101001011010010101011010,
64'b1001011001101001011010011001011001011010010110100101101001011010,
64'b0110011001100110011001100110011011110000111100001111000011110000,
64'b0110100101101001100101101001011010101010010101010101010110101010,
64'b0101010110101010010101011010101001011010101001011010010101011010,
64'b1001100101100110100110010110011001100110100110011001100101100110,
64'b0110011010011001100110010110011011111111000000001111111100000000,
64'b0011110000111100001111000011110001101001100101100110100110010110,
64'b0110011010011001100110010110011001100110011001100110011001100110,
64'b1100001111000011001111000011110010101010010101010101010110101010,
64'b0110011001100110011001100110011010011001100110010110011001100110,
64'b0101101010100101101001010101101000110011001100111100110011001100,
64'b1111000000001111000011111111000000000000000000000000000000000000,
64'b0011110011000011110000110011110011001100001100110011001111001100,
64'b0011110011000011110000110011110010011001011001101001100101100110,
64'b1001011010010110100101101001011011111111000000001111111100000000,
64'b0101101010100101101001010101101001011010101001011010010101011010,
64'b1100110011001100110011001100110000110011001100111100110011001100,
64'b1001100101100110100110010110011010101010010101010101010110101010,
64'b0011110011000011110000110011110011111111000000001111111100000000,
64'b0110100101101001100101101001011001010101010101011010101010101010,
64'b0101101010100101101001010101101001100110011001100110011001100110,
64'b0011110000111100001111000011110010100101101001010101101001011010,
64'b1111000000001111000011111111000001100110011001100110011001100110,
64'b1100110000110011001100111100110000001111111100000000111111110000,
64'b1010010101011010101001010101101000111100001111000011110000111100,
64'b0110011010011001100110010110011011110000000011110000111111110000,
64'b1010010110100101010110100101101011000011110000110011110000111100,
64'b1010101010101010101010101010101010100101010110101010010101011010,
64'b1001011010010110100101101001011001100110100110011001100101100110,
64'b1001011010010110100101101001011001011010010110100101101001011010,
64'b0101101010100101101001010101101010011001100110010110011001100110,
64'b1100110011001100110011001100110001010101010101011010101010101010,
64'b0000000011111111111111110000000011001100110011001100110011001100,
64'b0011110000111100001111000011110010010110100101101001011010010110,
64'b1001100101100110100110010110011000110011110011000011001111001100,
64'b1111000011110000111100001111000010010110100101101001011010010110,
64'b0110100110010110011010011001011000000000111111111111111100000000,
64'b1100001111000011001111000011110000001111111100000000111111110000,
64'b1010010101011010101001010101101000000000111111111111111100000000,
64'b0011110011000011110000110011110010100101010110101010010101011010,
64'b1100110011001100110011001100110010011001011001101001100101100110,
64'b1001100110011001011001100110011001101001011010011001011010010110,
64'b0000111111110000000011111111000010011001011001101001100101100110,
64'b0101010101010101101010101010101000111100001111000011110000111100,
64'b0110011010011001100110010110011001100110011001100110011001100110,
64'b1001011010010110100101101001011001011010010110100101101001011010,
64'b1111111111111111000000000000000011000011001111001100001100111100,
64'b1111111111111111000000000000000000001111000011111111000011110000,
64'b0000111100001111111100001111000011000011001111001100001100111100,
64'b1111000011110000111100001111000011111111111111110000000000000000,
64'b1010101010101010101010101010101010101010010101010101010110101010,
64'b0000000000000000000000000000000011111111111111110000000000000000,
64'b0101010110101010010101011010101001100110100110011001100101100110,
64'b1111000011110000111100001111000000111100001111000011110000111100,
64'b0011110000111100001111000011110001101001100101100110100110010110,
64'b1010101001010101010101011010101001101001011010011001011010010110,
64'b1100110011001100110011001100110000001111111100000000111111110000,
64'b0110100101101001100101101001011000111100001111000011110000111100,
64'b0110100110010110011010011001011000110011110011000011001111001100,
64'b0000000000000000000000000000000011110000000011110000111111110000,
64'b1010101010101010101010101010101011111111000000001111111100000000,
64'b0101010110101010010101011010101001011010101001011010010101011010,
64'b0101010110101010010101011010101000000000000000000000000000000000,
64'b1100110011001100110011001100110010011001100110010110011001100110,
64'b0000000000000000000000000000000010101010101010101010101010101010,
64'b0011001100110011110011001100110001101001011010011001011010010110,
64'b1111111100000000111111110000000010100101010110101010010101011010,
64'b0101010101010101101010101010101010010110011010010110100110010110,
64'b1111111111111111000000000000000011000011001111001100001100111100,
64'b1100001100111100110000110011110010101010010101010101010110101010,
64'b1111111111111111000000000000000000001111111100000000111111110000,
64'b1111111100000000111111110000000000001111000011111111000011110000,
64'b0101101010100101101001010101101000000000111111111111111100000000,
64'b1111000011110000111100001111000001010101010101011010101010101010,
64'b1100001100111100110000110011110011001100001100110011001111001100,
64'b1111111100000000111111110000000010101010101010101010101010101010,
64'b0101010110101010010101011010101000111100001111000011110000111100,
64'b0110011010011001100110010110011001100110011001100110011001100110,
64'b0101010101010101101010101010101011000011001111001100001100111100,
64'b0000000000000000000000000000000010011001011001101001100101100110,
64'b0011110011000011110000110011110000111100110000111100001100111100,
64'b0110011001100110011001100110011001011010101001011010010101011010,
64'b1100001111000011001111000011110000110011001100111100110011001100,
64'b0011110011000011110000110011110010101010010101010101010110101010,
64'b0011110000111100001111000011110011111111000000001111111100000000,
64'b1001011010010110100101101001011001010101010101011010101010101010,
64'b0110100110010110011010011001011001100110011001100110011001100110,
64'b0000000000000000000000000000000010100101101001010101101001011010,
64'b0011001111001100001100111100110001100110011001100110011001100110,
64'b1001011001101001011010011001011000001111111100000000111111110000,
64'b1010010101011010101001010101101000111100001111000011110000111100,
64'b1100001111000011001111000011110011110000000011110000111111110000,
64'b0000000000000000000000000000000000111100001111000011110000111100,
64'b0101101010100101101001010101101000000000000000000000000000000000,
64'b1001011010010110100101101001011010101010010101010101010110101010,
64'b0000111111110000000011111111000011000011001111001100001100111100,
64'b0101101010100101101001010101101010100101010110101010010101011010,
64'b1010010101011010101001010101101000111100001111000011110000111100,
64'b1100001100111100110000110011110010010110011010010110100110010110,
64'b0011110011000011110000110011110010101010101010101010101010101010,
64'b0000000000000000000000000000000011000011110000110011110000111100,
64'b0000111100001111111100001111000001011010101001011010010101011010,
64'b0011110011000011110000110011110010100101101001010101101001011010,
64'b0110011010011001100110010110011001101001011010011001011010010110,
64'b0000111111110000000011111111000010100101010110101010010101011010,
64'b1010101010101010101010101010101000001111111100000000111111110000,
64'b1001011010010110100101101001011001011010101001011010010101011010,
64'b1010010101011010101001010101101011111111111111110000000000000000,
64'b1001100110011001011001100110011011000011110000110011110000111100,
64'b1111000011110000111100001111000011110000111100001111000011110000,
64'b0000111111110000000011111111000001100110100110011001100101100110,
64'b1010101010101010101010101010101001100110011001100110011001100110,
64'b1100110000110011001100111100110001011010010110100101101001011010,
64'b0101101010100101101001010101101011111111111111110000000000000000,
64'b0011001100110011110011001100110010101010101010101010101010101010,
64'b1111111111111111000000000000000000111100001111000011110000111100,
64'b0000111111110000000011111111000000001111000011111111000011110000,
64'b0000111111110000000011111111000011000011001111001100001100111100,
64'b0110011001100110011001100110011001010101101010100101010110101010,
64'b1001100110011001011001100110011001100110100110011001100101100110,
64'b0000000011111111111111110000000010101010101010101010101010101010,
64'b1010010101011010101001010101101010100101010110101010010101011010,
64'b0110100101101001100101101001011001010101101010100101010110101010,
64'b0110100110010110011010011001011011000011110000110011110000111100,
64'b1001011001101001011010011001011010010110100101101001011010010110,
64'b0011001100110011110011001100110000110011110011000011001111001100,
64'b1001011010010110100101101001011000000000000000000000000000000000,
64'b1001011001101001011010011001011001100110011001100110011001100110,
64'b0000111111110000000011111111000000001111111100000000111111110000,
64'b1100110011001100110011001100110011111111000000001111111100000000,
64'b1010010101011010101001010101101001011010101001011010010101011010,
64'b1001011010010110100101101001011011001100110011001100110011001100,
64'b0011110000111100001111000011110011000011110000110011110000111100,
64'b0101010101010101101010101010101001100110011001100110011001100110,
64'b0110011010011001100110010110011011001100001100110011001111001100,
64'b1100001100111100110000110011110000110011001100111100110011001100,
64'b1001011001101001011010011001011000001111111100000000111111110000,
64'b0011110011000011110000110011110001101001100101100110100110010110,
64'b0101101001011010010110100101101000001111000011111111000011110000,
64'b0110100110010110011010011001011000000000000000000000000000000000,
64'b0011110011000011110000110011110000111100001111000011110000111100,
64'b1010101001010101010101011010101000000000111111111111111100000000,
64'b1111000011110000111100001111000011111111111111110000000000000000,
64'b1100110000110011001100111100110011001100001100110011001111001100,
64'b1100001100111100110000110011110001011010010110100101101001011010,
64'b0101010101010101101010101010101001010101010101011010101010101010,
64'b0000000000000000000000000000000001011010010110100101101001011010,
64'b1111000000001111000011111111000010010110011010010110100110010110,
64'b0110011001100110011001100110011001100110100110011001100101100110,
64'b0101010110101010010101011010101011000011001111001100001100111100,
64'b0000000000000000000000000000000001100110011001100110011001100110,
64'b1010010101011010101001010101101011000011001111001100001100111100,
64'b1100110011001100110011001100110001011010101001011010010101011010,
64'b0011110000111100001111000011110011000011110000110011110000111100,
64'b0011110011000011110000110011110001011010101001011010010101011010,
64'b0011001100110011110011001100110011001100001100110011001111001100,
64'b1010101010101010101010101010101000000000000000000000000000000000,
64'b0000111111110000000011111111000000110011110011000011001111001100,
64'b0011110011000011110000110011110011001100110011001100110011001100,
64'b0110011001100110011001100110011010011001011001101001100101100110,
64'b1001100110011001011001100110011000111100110000111100001100111100,
64'b1010101001010101010101011010101001101001011010011001011010010110,
64'b0101101001011010010110100101101001011010101001011010010101011010,
64'b0101101010100101101001010101101000111100001111000011110000111100,
64'b1111000000001111000011111111000011110000000011110000111111110000,
64'b0000000011111111111111110000000011001100001100110011001111001100,
64'b1100001111000011001111000011110010100101010110101010010101011010,
64'b0101010101010101101010101010101001100110100110011001100101100110,
64'b0011110011000011110000110011110010100101101001010101101001011010,
64'b1100001111000011001111000011110010101010101010101010101010101010,
64'b0101010110101010010101011010101011110000111100001111000011110000,
64'b0000000000000000000000000000000001011010010110100101101001011010,
64'b0101101001011010010110100101101011000011110000110011110000111100,
64'b1010010101011010101001010101101011110000000011110000111111110000,
64'b1010010101011010101001010101101001101001100101100110100110010110,
64'b1111000000001111000011111111000001100110100110011001100101100110,
64'b1001011010010110100101101001011010100101010110101010010101011010,
64'b1001011001101001011010011001011000000000111111111111111100000000,
64'b1010010101011010101001010101101010100101101001010101101001011010,
64'b0110100101101001100101101001011001100110100110011001100101100110,
64'b1100001100111100110000110011110011000011110000110011110000111100,
64'b0011110000111100001111000011110010011001011001101001100101100110,
64'b0000000011111111111111110000000001100110011001100110011001100110,
64'b1100110011001100110011001100110011111111000000001111111100000000,
64'b0000000000000000000000000000000010011001011001101001100101100110,
64'b0011001111001100001100111100110000001111111100000000111111110000,
64'b1100110000110011001100111100110010101010010101010101010110101010,
64'b1100110000110011001100111100110010010110011010010110100110010110,
64'b0000000011111111111111110000000011000011110000110011110000111100,
64'b0110100110010110011010011001011001100110100110011001100101100110,
64'b0011110011000011110000110011110011111111111111110000000000000000,
64'b0110011010011001100110010110011010011001011001101001100101100110,
64'b1100001100111100110000110011110001101001011010011001011010010110,
64'b0101101010100101101001010101101010100101010110101010010101011010,
64'b0000111111110000000011111111000001101001011010011001011010010110,
64'b1111111111111111000000000000000000111100001111000011110000111100,
64'b0101101001011010010110100101101000000000000000000000000000000000,
64'b0000000000000000000000000000000001101001011010011001011010010110,
64'b0000111100001111111100001111000000000000111111111111111100000000,
64'b0000111100001111111100001111000000110011001100111100110011001100,
64'b1010010110100101010110100101101010010110011010010110100110010110,
64'b0101010101010101101010101010101010100101010110101010010101011010,
64'b1001011001101001011010011001011001101001011010011001011010010110,
64'b1111000000001111000011111111000010101010101010101010101010101010,
64'b0110100101101001100101101001011001101001011010011001011010010110,
64'b0101101010100101101001010101101011000011001111001100001100111100,
64'b1100110000110011001100111100110001100110100110011001100101100110,
64'b1010101001010101010101011010101011000011001111001100001100111100,
64'b0000000000000000000000000000000010100101010110101010010101011010,
64'b1001100101100110100110010110011000000000000000000000000000000000,
64'b0000000000000000000000000000000011000011001111001100001100111100,
64'b1111111100000000111111110000000001010101010101011010101010101010,
64'b0101010110101010010101011010101001011010010110100101101001011010,
64'b1001100101100110100110010110011010010110011010010110100110010110,
64'b0110011001100110011001100110011001100110100110011001100101100110,
64'b1001011001101001011010011001011011000011001111001100001100111100,
64'b1010101001010101010101011010101001100110011001100110011001100110,
64'b0110100110010110011010011001011011000011001111001100001100111100,
64'b0110011010011001100110010110011001011010101001011010010101011010,
64'b1010010110100101010110100101101011000011110000110011110000111100,
64'b1001100110011001011001100110011001011010101001011010010101011010,
64'b1010101010101010101010101010101011001100001100110011001111001100,
64'b0011110000111100001111000011110000000000000000000000000000000000

} ;
























parameter  [0:SEG_NUM*32-1] D_CRC_REG_INIT = { 

32'b01101001000001001011101101011001,
32'b01010101001011010010001011001000,
32'b11111011101011000111110000111010,
32'b01001010010101011010111101100111,
32'b01110010010000111100100001101000,
32'b01010110001100101110111010110000,
32'b01101101010110101110110000110100,
32'b10010011001110010100111001010001,
32'b10110101001000101011110000001111,
32'b10011000111001110011101110001110,
32'b01001101111001011011110100100000,
32'b10001010010110011101000010100010,
32'b00001011101111110000011100010100,
32'b01000010010010101000001000100111,
32'b00011011101000010100010101100011,
32'b01000110101000001110101010111100,
32'b10011000001100110011001100010001,
32'b11000110010111111010111111110001,
32'b01100100101101101100000100010111,
32'b00111001001101010001111110101010,
32'b11010110110000110110100010001111,
32'b00001001100001011111010100001011,
32'b10010010000011011100011111110101,
32'b10110000111011110000000000101110,
32'b10010001111010100111000101101100,
32'b01100010100011101011101100000101,
32'b01001001000000010101011011011110,
32'b00111001001001010111101101000011,
32'b11100100000010010101010000001110,
32'b00110111110110110111100111000010,
32'b11011100010011000010000110100010,
32'b11100101010111101001011001001111,
32'b11111010001111001111100110101111,
32'b11101111101010101000010011110001,
32'b11001001010101001010000011011110,
32'b10110101101010011011000000101000,
32'b01011010100100010110001010100101,
32'b00011101100111010111010100011101,
32'b01010100001011111111101011001101,
32'b01001101000101010001110001001010,
32'b00011101101010101011011001010010,
32'b01110110111010101110101101001011,
32'b01111000101001101011100011111011,
32'b01101001100111010100101000100000,
32'b10011100000111010010001100010111,
32'b10110100100110011010001111011000,
32'b00111111101101100110110001110010,
32'b00011101011101001010001011101110,
32'b11001011000101000110111101110001,
32'b11001111010011111011101110011101,
32'b10110011101110100100111010001100,
32'b10110110111001110101000010011110,
32'b11010100001100010000110100011011,
32'b11010110100110111010011100010010,
32'b01000011110001100000101110111001,
32'b00111101100101111010111010011101,
32'b11011100011010111001101010001010,
32'b00001000011000110110001001111100,
32'b00110000001011100110011000101000,
32'b01001110001111001010001000100000,
32'b00101011001001101100010111010100,
32'b10100010101101101110110000101011,
32'b00000100111100000110100001110111,
32'b11100001010100011010101010110010

 } ;




































parameter [0:GO_BACK_STAGE*256*64-1] GO_BACK_POLY_STRIDE_8 = 
{
    
64'b0000000001101100011010100000101000001100011011001100000001100000,
64'b0110110010100000011001101010000000001010101011001010101010100000,
64'b1100101010100000011000001100000001101010011011001010110010100000,
64'b1010000001100000110010100000000000001100101010100000101011000000,
64'b1100101011000000101001101010000010100000011010100110101000000000,
64'b1100000011000000000001100110000001101010011010101010000001100000,
64'b1100011000001100011001101100000000000110110000001010011001100000,
64'b1010110001101100101010100000000011000110011010101100110011000000,
64'b0110000001101100011000001100000000001010101001101010000010101010,
64'b1010011011000000011011000000000001101010000010100000110001100000,
64'b1010101001100000110001100110000010100110110001101100101011000000,
64'b1100000000000000011010100110000010100110110000000000101000000000,
64'b0110000010101100011011000000000000000110000011000110011000000000,
64'b1100110011001100011001100110000010100000000011000110110010100000,
64'b1010011001100000000001101100000000000110011000001010101010100000,
64'b0000110000000110000000001100000010100110000001101010000001100000,
64'b1010000000001100101011001010110010101010011010101010000001100000,
64'b1010110011001010000010100110000000000110011010100110110001100000,
64'b0110110001100000000010101100000011001100110010101100000011000000,
64'b1100000010100000011001101010000010100000011001100000011000000000,
64'b1100011001100000110010100110000011001010110011001100110010100000,
64'b0110000001100000000000001010000011001100011011000110000011000000,
64'b0110101010101100101000000110000010101100101000001100110001100000,
64'b1100011010100110110011001010000000000110011011000000101010100000,
64'b1010101000000110101000001100000010100110011011000110101001101100,
64'b1100101001101010000011001010000011001100000001100000000011000000,
64'b0110110000000000011000001010000001101100000011000000011010100000,
64'b1100000010100000000011000000000011000110101010101010110010100000,
64'b0000000001101100000011001010000000000110101000001100110000000000,
64'b0110110011000110000000001010000011001010000010100110101011000000,
64'b1100000000001010101000000110000000001100110010100110011011000000,
64'b0000011010101010000010100110000011000110101011001100000011000000,
64'b1100101001100110101010101100000011001100110011001100000011000000,
64'b1010110010100110011000000110101000001100011011001100000001100000,
64'b0000000011000000011011000110000000001010101011001010101010100000,
64'b0000101000000000000001100110000001101010011011001010110010100000,
64'b0110011000000000000000000110000000001100101010100000101011000000,
64'b1010101010100000101001100000000010100000011010100110101000000000,
64'b1010101001101100101001100000000001101010011010101010000001100000,
64'b0000000010101010101010100110000000000110110000001010011001100000,
64'b0000011001101010000010101100000011000110011010101100110011000000,
64'b1010101000000110011011000110000000001010101001101010000010101010,
64'b1100101011000000000011001010000001101010000010100000110001100000,
64'b0110101011000000110010100110000010100110110001101100101011000000,
64'b1100000001101100011001101100000010100110110000000000101000000000,
64'b0000110001101010011011001010000000000110000011000110011000000000,
64'b0000110011000110110001100000000010100000000011000110110010100000,
64'b1010000011001010000011001010000000000110011000001010101010100000,
64'b0000110011001100011001101010000000001010000010100000000010100000,
64'b0110000001100110110000000110110010101010011010101010000001100000,
64'b0000101000001010011000000110000000000110011010100110110001100000,
64'b0000110010100000101001100110000011001100110010101100000011000000,
64'b1100110000000000000010100110000010100000011001100000011000000000,
64'b0110011011000000110011001010000011001010110011001100110010100000,
64'b1100110011000000110001100000000011001100011011000110000011000000,
64'b0000000001100110110001101100000010101100101000001100110001100000,
64'b0000110011001100000011001010000000000110011011000000101010100000,
64'b1100011010101100110000000110000010100110011011000110101001101100,
64'b0000110000001010101010100110000011001100000001100000000011000000,
64'b0110110010100000000001101100000001101100000011000000011010100000,
64'b1010000001100000011011001010000011000110101010101010110010100000,
64'b1010000001100110011010100110000000000110101000001100110000000000,
64'b0000101010101100101001100000000011001010000010100110101011000000,
64'b1100101010100110101010101100000000001100110010100110011011000000,
64'b0000101011000110101001101100000010101100000011001010000001100000,
64'b1010011011000110110011000110000011001100110011001100000011000000,
64'b0110011000000110000000001010101000001100011011001100000001100000,
64'b1010000010100000101001100110000000001010101011001010101010100000,
64'b1100000011000000101000001100000001101010011011001010110010100000,
64'b1010011011000000000001100000000000001100101010100000101011000000,
64'b0110110010101100110000001100000010100000011010100110101000000000,
64'b0000011000000000000011000000000001101010011010101010000001100000,
64'b0110000011000110110010101010000000000110110000001010011001100000,
64'b1010000010101010011001101100000011000110011010101100110011000000,
64'b0000000001100110101010100000000000001010101001101010000010101010,
64'b0000101011000000011001101100000001101010000010100000110001100000,
64'b0000101001101100101001100110000010100110110001101100101011000000,
64'b0000110010100000000000001010000010100110110000000000101000000000,
64'b1010101000001010011010100110000000000110000011000110011000000000,
64'b0000000011000000110001101100000010100000000011000110110010100000,
64'b0000011001100000000011000000000001100000101010100110000001100000,
64'b1010000000000110011011001100000000001010000010100000000010100000,
64'b0000110000000110110010101010110010101010011010101010000001100000,
64'b1100101010101010000001101100000000000110011010100110110001100000,
64'b1100101011000000011011000000000011001100110010101100000011000000,
64'b1010110001100000000010101100000010100000011001100000011000000000,
64'b0000110001101100011011001100000011001010110011001100110010100000,
64'b0000101001100110000010101010000011001100011011000110000011000000,
64'b1010101001100000011001100000000010101100101000001100110001100000,
64'b1100011010100110000000000000000000000110011011000000101010100000,
64'b1010101010101100101000001100000010100110011011000110101001101100,
64'b1100110010101010101001100110000011001100000001100000000011000000,
64'b0110110011001100000010100110000001101100000011000000011010100000,
64'b1100110010100110011011000000000011000110101010101010110010100000,
64'b0110000001101100110010100000000000000110101000001100110000000000,
64'b0000110000000110101011000110000011001010000010100110101011000000,
64'b0000110001100000101010100000000011001010000010100000101001100000,
64'b1100101010101100110010100000000011000000101011001100011011000000,
64'b0000000000000110101001100110000000000110011011001010000000000000,
64'b0000011011000110101011000000101010101100000011000000101001100000,
64'b1010110000000000110010101010000011000000011011000000110000000000,
64'b0110000001100000101001100000000010101010101011001010101011000000,
64'b0000101001100000110000001010000011001010101001100110110000000000,
64'b0000011001100110101001100110000000001100000001101100000000000000,
64'b1100110001101010110011000000000000001010000001101100000010100000,
64'b0000110001101100101010100000000010100000000000001100101001100000,
64'b0110011011001010110000000000000001101100000010100000101010100000,
64'b0000000011000110110011000110000011001010101001101100101011001010,
64'b0110101000000000000001100110000000001010101001100110000001100000,
64'b1010101001100110110000001010000001101010000010101010110010100000,
64'b0110101011001010101001100000000000000000101000000000110011000000,
64'b1010000010100110011000001100000000001010000010100110011011000000,
64'b1010000000000110101011001010000000000110011000000110110011000000,
64'b0110101011000000011010101010000011001100011000000110101000000000,
64'b0110101010100110000011000000000001100110011010100000101001100000,
64'b1010110001100110000000001010110001101010110010101100011011000000,
64'b0000000001101010101000000110000011000000000010101010011000000000,
64'b0000101000000000011010100110000010101100101010101100000001100000,
64'b0110101001101100011011000000000011001010110010101010011001100000,
64'b1010000000000000110001101100000000001100011010100000000000000000,
64'b0110101000001010011010100110000001100110011010101100000000000000,
64'b0000110010100000000010100000000001100110110010101100000011000000,
64'b0110110011000110110001100110000001101010011011000110101000000000,
64'b0110101010101100110010101010000001100110110011000110011001101100,
64'b1010110000000110110010100110000011001100011010100000110001100000,
64'b1010000000000000011011000000000000000000110010100000011000000000,
64'b0110101011000110011010101100000000000110101000000000110011000000,
64'b0110110001101010110010101100000000000000000010101100011001100000,
64'b0110101001101010101000001100000010100110011000001100000000000000,
64'b1010000010101010101000000110000000001010011000000110011010100000,
64'b1010011011001100110000001100000001100110011011001010110011000000,
64'b1100000010100110110000001100000001100110101011000000110010100000,
64'b1100000010100110011001100110101010100000101011000110011010100000,
64'b1100110001100000110010100000000001100000110011000000101011000000,
64'b0000101011001100000001100110000000000110000011000110110001100000,
64'b1100110011000110000011000000000010100000011011000000101010100000,
64'b1010110001100000000001101010000011000110011011000000000000000000,
64'b0000011000000000110000001010000001100110101011001010000000000000,
64'b0110000001101100110010101010000001100110011000000110110010100000,
64'b1010011001101010110011000000000001101100101010100110110011000000,
64'b0000000010101010110000001100000010101010011001101010101001101010,
64'b0000011011000110000001101100000010101010101011000000011010100000,
64'b0110101001101100011000001100000000001100011000000000101000000000,
64'b0110110001100000101011000110000000001010000011000000011001100000,
64'b1100110001100110110000000000000011001100110010100000000000000000,
64'b0110000001101100110000000110000000000110011000000110110011000000,
64'b1100110000000000000000001010000011001100011000000110101000000000,
64'b0000101001100110101000001010000001100110011010100000101001100000,
64'b1010000011000110011011000110110001101010110010101100011011000000,
64'b1010000011001010101001101010000011000000000010101010011000000000,
64'b1010011010100000101011001100000010101100101010101100000001100000,
64'b0000000010100110000010101010000011001010110010101010011001100000,
64'b0110101001101010000001101100000000001100011010100000000000000000,
64'b0000011010100000000010101100000001100110011010101100000000000000,
64'b1100101011000000101011001100000001100110110010101100000011000000,
64'b0110110001100110101000000000000001101010011011000110101000000000,
64'b0000101001101100101010100000000001100110110011000110011001101100,
64'b0000110000001100101011001010000011001100011010100000110001100000,
64'b1100011001101010110010101010000000000000110010100000011000000000,
64'b0110000001101010011000000110000000000110101000000000110011000000,
64'b0000000000000000110010101010000010100000011000001100101000000000,
64'b0000011011001010110001100110000011001010110000001010011010100000,
64'b0110101000001010110000001010000011000000110000000000011001100000,
64'b0000011010101100000010101100000011000110000011000110011011000000,
64'b0000101001100110011001100110000010101100011011001010101000000000,
64'b0000000001100110011000000000101001100000011011000110000011000000,
64'b0000101001101100101011001100000010100110110000000110110000000000,
64'b1010011010100000101011000110000010101010011000001100011001100000,
64'b1010110010101010011011001100000011000000000000000110101001100000,
64'b0000101010100000011010101010000001100000101011000110110000000000,
64'b1010110001100000000001101100000011001100110011000110011001100000,
64'b1010000001101100101000001100000010100110011000000000011011000000,
64'b1100011011000110101000000000000000001100000001100000000011000000,
64'b1100110001100110101001101010000001100110101010101100110000001010,
64'b1010000010100110000000000000000000001100110011000000000001100000,
64'b0110011001101010011000000000000000000000011001100000101011000000,
64'b0000000011001100110001100110000001100000110000001010110010100000,
64'b0110000010101100110010100110000000001100101000000110110011000000,
64'b0000110000001100110010101010000010100000101000000000011011000000,
64'b0000110010100000011001100000000010101100101000001100011010100000,
64'b1100110000000110011010101100000001101010110010100110011010100000,
64'b1100000010100110011011001100110011001010011010101100000000000000,
64'b1100101001100110000001101100000001101100101010100110000010100000,
64'b0110000000000110011000000110000011000110011000001010011011000000,
64'b1010101010100000101010100110000000000000101000000110011001100000,
64'b1010000000000000000010100110000001100000110000000110000010100000,
64'b0110101010100000011010100110000010100000000010100110011011000000,
64'b0000101001100000101000001100000001100110011010101010011010100000,
64'b0110110000001010101011001010000000001010101011000000101010100000,
64'b0110011010101010101010101010000011000110110001100000000010101100,
64'b1100110000000110000011001100000010101010000000001010101011000000,
64'b1100000011000000110000001100000000001010011001100000110010100000,
64'b1010000011001100110011000110000011001010101000000110000011000000,
64'b1010110011001010110000001100000010100000011000001100101000000000,
64'b0110101010101010110011001010000011001010110000001010011010100000,
64'b1010101010101010101001100000000011000000110000000000011001100000,
64'b1100000011001100110000001010000011000110000011000110011011000000,
64'b0110101000000110011001101100000010101100011011001010101000000000,
64'b0110101011001010110000000110101001100000011011000110000011000000,
64'b1100110011001010011000000110000010100110110000000110110000000000,
64'b0000110010100110000011001010000010101010011000001100011001100000,
64'b0110011011000000011000000110000011000000000000000110101001100000,
64'b0110011010100000000010100000000001100000101011000110110000000000,
64'b0110110011000000000010101100000011001100110011000110011001100000,
64'b1010000000000000101011000110000010100110011000000000011011000000,
64'b1010101000000000101000001010000000001100000001100000000011000000,
64'b0000110001101100000001101100000001100110101010101100110000001010,
64'b1010011000001100000010100110000000001100110011000000000001100000,
64'b0110101000001010101010101100000010100110110000000110101000000000,
64'b1100000010100110101010101010000001100000110000001010110010100000,
64'b1100011001101100101000000110000000001100101000000110110011000000,
64'b0110110011001100011001100000000010100000101000000000011011000000,
64'b0000000000000000000010101100000010101100101000001100011010100000,
64'b0110110010100110011011000000000001101010110010100110011010100000,
64'b0110110000000110101010100110110011001010011010101100000000000000,
64'b1010000010101100011000000110000001101100101010100110000010100000,
64'b1010101001101100101000000110000011000110011000001010011011000000,
64'b1100011000001010110010101100000000000000101000000110011001100000,
64'b0110011001100000101011001010000001100000110000000110000010100000,
64'b0110101000000000000011000000000010100000000010100110011011000000,
64'b0110101010100000110000000110000001100110011010101010011010100000,
64'b1100110000000000110010100110000000001010101011000000101010100000,
64'b0000000011000000000011000000000011000110110001100000000010101100,
64'b1100011010101010000001100110000010101010000000001010101011000000,
64'b0110011000001100110011000000000001101100101000000110011010100000,
64'b1010000011001100110011000110000011001010101000000110000011000000,
64'b1010110011001010110000001100000010100000011000001100101000000000,
64'b0110101010101010110011001010000011001010110000001010011010100000,
64'b1010101010101010101001100000000011000000110000000000011001100000,
64'b1100000011001100110000001010000011000110000011000110011011000000,
64'b0110101000000110011001101100000010101100011011001010101000000000,
64'b0110101011001010110000000110101001100000011011000110000011000000,
64'b1100110011001010011000000110000010100110110000000110110000000000,
64'b0000110010100110000011001010000010101010011000001100011001100000,
64'b0110011011000000011000000110000011000000000000000110101001100000,
64'b0110011010100000000010100000000001100000101011000110110000000000,
64'b0110110011000000000010101100000011001100110011000110011001100000,
64'b1010000000000000101011000110000010100110011000000000011011000000,
64'b1010101000000000101000001010000000001100000001100000000011000000,
64'b0000110001101100000001101100000001100110101010101100110000001010,
64'b1100011000000000000000001010000011000000011010100110110011000000,
64'b0110101000001010101010101100000010100110110000000110101000000000,
64'b1100000010100110101010101010000001100000110000001010110010100000,
64'b1100011001101100101000000110000000001100101000000110110011000000,
64'b0110110011001100011001100000000010100000101000000000011011000000,
64'b0000000000000000000010101100000010101100101000001100011010100000,
64'b0110110010100110011011000000000001101010110010100110011010100000,
64'b0110110000000110101010100110110011001010011010101100000000000000,
64'b1010000010101100011000000110000001101100101010100110000010100000,
64'b1010101001101100101000000110000011000110011000001010011011000000,
64'b1100011000001010110010101100000000000000101000000110011001100000,
64'b0110011001100000101011001010000001100000110000000110000010100000,
64'b0110101000000000000011000000000010100000000010100110011011000000,
64'b0110101010100000110000000110000001100110011010101010011010100000,
64'b1100110000000000110010100110000000001010101011000000101010100000,
64'b0000000011000000000011000000000011000110110001100000000010101100,
64'b1010011001100110110011001100101010101100000000001100101010100000,
64'b0000000010101100011000001010000011000110000011000110110000000000,
64'b1100000011000110000010101010000011000000110011000110011000000000,
64'b1100110001100110011000001100000010101100101010100000110011000000,
64'b0000000011001100101000001010000000000000000010100110000000000000,
64'b1010110001100000110001101100000010100110110011000110110000000000,
64'b1010110001101100000010100110000000001010101000001010011000000000,
64'b0000110000000000011010101010000001100000110000000000000000000000,
64'b0110011010101100000011001100000011001010101001101010101001101010,
64'b1010101011000110110010101100000011001010101010100110101011000000,
64'b1010101011001100011011000000000000001100110011000000000010100000,
64'b0110110011000000110001100000000011000000000001100110000011000000,
64'b0110000000001100011000000110000011000110110000001010011010100000,
64'b0000110010101010000010100110000011000110011000000110101001100000,
64'b0000000000001100110010100110000010101010011010101010110010100000,
64'b0110101010101010101010100110000011000000101000000110000000000000,
64'b0110000010100000110011001100110001101010101010100000110011000000,
64'b0000101011000110000010101100000000000110000000000110000000000000,
64'b1100000011000000101001100110000010101010000010100110011000000000,
64'b0110110000000000101000001100000001100000011001101010101000000000,
64'b1010101001100110110000001100000000001010000011001100101010100000,
64'b0110110000001010110010101100000011001100000000000110000000000000,
64'b0110011000001100101011000000000000000110011010100110011000000000,
64'b0000011010101010101001101100000011000000000000000000101000000000,
64'b1010000001101100101011001100000010101100011011001100110011001100,
64'b1100110011000000110011000110000010101100110001101100110010100000,
64'b0110011001100110000011001010000010100000000000001010000001100000,
64'b1010110001101010011000000000000000001010101001101100000000000000,
64'b0000101010101100000010101010000010101100000010100110110001100000,
64'b1010110001101100101001100000000010100110011000001100011011000000,
64'b0000101000001100110001100000000001100110011011000110000001100000,
64'b1010011001101100110001100000000000000000011000001100101000000000,
64'b0110110010101100011011000110000001101100011011000000000010100000,
64'b1010110010100000110001100000101010101100000000001100101010100000,
64'b1100000001101100110001101100000011000110000011000110110000000000,
64'b1010110011000110101010100110000011000000110011000110011000000000,
64'b0110011000000000101000000000000010101100101010100000110011000000,
64'b0110110011000110011010100110000000000000000010100110000000000000,
64'b1100101001101100011010101100000010100110110011000110110000000000,
64'b1010101011000110101011001010000000001010101000001010011000000000,
64'b1010110001101100110001100110000001100000110000000000000000000000,
64'b1010101001101100110000001010000011001010101001101010101001101010,
64'b1100110010100000110001100110000011001010101010100110101011000000,
64'b0000011010100110000011000000000000001100110011000000000010100000,
64'b0110011001101100110011001010000011000000000001100110000011000000,
64'b1100110001100000110001100110000011000110110000001010011010100000,
64'b0000011010100110110011000110000011000110011000000110101001100000,
64'b1010011001100000000011000110000010101010011010101010110010100000,
64'b1100101011000000110010101100000001100000110000000000101001100000,
64'b0110101011001010101001101010110001101010101010100000110011000000,
64'b0000101011000000101001100000000000000110000000000110000000000000,
64'b0110000010100110011001100110000010101010000010100110011000000000,
64'b1100011010101010110000001010000001100000011001101010101000000000,
64'b0110101000001100110011001100000000001010000011001100101010100000,
64'b1010011001101010011011001010000011001100000000000110000000000000,
64'b0110110010100110011000000110000000000110011010100110011000000000,
64'b1100000001101010000001101100000011000000000000000000101000000000,
64'b1100011001101010101010100110000010101100011011001100110011001100,
64'b0000000001101010101011001100000010101100110001101100110010100000,
64'b1010011011001100101010101010000010100000000000001010000001100000,
64'b1100011011001010000010101100000000001010101001101100000000000000,
64'b1010101001101010101001101100000010101100000010100110110001100000,
64'b1010011001101100101010100110000010100110011000001100011011000000,
64'b1100011011001010101010100110000001100110011011000110000001100000,
64'b0000101001100110110000000110000001100000101000001010011011000000,
64'b0110110000000000000011001100000001101100011011000000000010100000,
64'b0110110001100110110011001010101010101100000000001100101010100000,
64'b0000110000001010101001100000000011000110000011000110110000000000,
64'b1010110000001010000010101100000011000000110011000110011000000000,
64'b1100101001100000011001101100000010101100101010100000110011000000,
64'b1100000010101010011000000000000000000000000010100110000000000000,
64'b1100011001101100000000000110000010100110110011000110110000000000,
64'b1100110001101010101000000110000000001010101000001010011000000000,
64'b0000011010101010000011001010000001100000110000000000000000000000,
64'b0000000010100000101011001010000011001010101001101010101001101010,
64'b1010000001100000000000000110000011001010101010100110101011000000,
64'b0110011010101010011011000110000000001100110011000000000010100000,
64'b0110101011000110110001101100000011000000000001100110000011000000,
64'b1100110001101100000011000000000011000110110000001010011010100000,
64'b0110110000001100011001100000000011000110011000000110101001100000,
64'b0000101000001010110011001010000001100000110000000110110010100000,
64'b1100000000000110110000000000000001100000110000000000101001100000,
64'b1010101000001010000000001100110001101010101010100000110011000000,
64'b0110011011000000000001101100000000000110000000000110000000000000,
64'b1100101011000000101001101010000010101010000010100110011000000000,
64'b1010101010100000000010100110000001100000011001101010101000000000,
64'b0000110000000000011000001100000000001010000011001100101010100000,
64'b1010000011000000110010100110000011001100000000000110000000000000,
64'b1100110011001010110011001010000000000110011010100110011000000000,
64'b0000110010101010110010101010000011000000000000000000101000000000,
64'b1010000000001100101001101100000010101100011011001100110011001100,
64'b1010110000000000110011001100000010101100110001101100110010100000,
64'b1010110001100000101000000000000010100000000000001010000001100000,
64'b0110101010100110101011001100000000001010101001101100000000000000,
64'b1010000001100110011000001100000010101100000010100110110001100000,
64'b0000000000000000011011000110000010100110011000001100011011000000,
64'b1010110010101100000010100110000001100110110011001010011000000000,
64'b0000000000001100101010100000000001100000000011001100011001100000,
64'b0110110000000110101000000000000010101100101010100000101000000000,
64'b1100110000000000000011001010101001100000011001101010101001100000,
64'b1010011010100000110001100110000011000110110000001100110010100000,
64'b0110110001100000000001101100000001101100101011001010000011000000,
64'b0000000000000000110000001010000000000000110001100000011010100000,
64'b1100101000000000101011000110000000001100000010100000101010100000,
64'b0000000010101100101000000110000011000000011000000110000011000000,
64'b1010101001101100101001101100000010100000011001100110110011000000,
64'b1100101000000000011011000000000011001010000011000110110000000000,
64'b1100000000001010000010101010000010100110011001100110110001101010,
64'b1100101011000000011010101010000010101010101001100000101010100000,
64'b1100011001101100110000000000000000000000011001100000101011000000,
64'b0110000011000110110010101010000011000000000010101010101010100000,
64'b0000000010101010011000000110000010101100011010100000110011000000,
64'b0110011010100110011000000000000011000000011011001010000011000000,
64'b0000101010100110101011000000000001101010000001100110011001100000,
64'b0000000011000000110010101010000010100000000000001010110000000000,
64'b0110011001101100011000000000110000000110101010101010110000000000,
64'b0110011000001100101001100110000010101100011001101010000011000000,
64'b0110011010100000011000000110000011000110000000001010110011000000,
64'b0000011011001100000000000000000000000110011010100000011000000000,
64'b0000000000000000000010100110000000001100101001100110110001100000,
64'b1100011001101100110001101010000001101100011011001100110011000000,
64'b0110011000001100000001100110000011001010101010101010101001100000,
64'b1010011001100110101001101010000010100110011001100000011010100000,
64'b1100110011001100011000001100000000000000000001101010110011001100,
64'b1100110000001100101011001010000010100110011010101100011000000000,
64'b1010000011001010101010100110000000001100011011000000011001100000,
64'b0110101010101010011001101010000000000000101010100000011000000000,
64'b1100101011001100110010101010000000001010011001101010101001100000,
64'b1100000010101010000001100110000000000000011000001100000000000000,
64'b1010011001101010000000001010000001101100101001101100110001100000,
64'b1100000011001100000011000110000001100000000010100110101010100000,
64'b0000000000000110000000001100000000001100110011001100101000000000,
64'b0110011001100110110011000110101011001010110011001100101000000000,
64'b1100101010101010000011001010000000000110101010101100000010100000,
64'b0000101001101100101010101100000010100110110011000000011010100000,
64'b0000011010101010011001100110000000001010011011001100101011000000,
64'b0110101001101100000000001010000011001010110010101010101010100000,
64'b1100110001101100011011000000000010100110011001100110011001100000,
64'b1100110000001010101010100110000001101100110011000000110001100000,
64'b0110011001101010000011000000000000001010101001101100101000000000,
64'b1100101010100110000000000000000011001100110001100000011010101010,
64'b0110011010101100110011001010000000001010011000001010011011000000,
64'b1100110001100000000001100000000000001010011001100000011010100000,
64'b1100011010101010000011001010000000001100110011001100011011000000,
64'b1010101001100110000011001100000010100000110000000000101000000000,
64'b0110110011001100000010100110000011000000011011001010000011000000,
64'b0000101010100000000000001100000001101010000001100110011001100000,
64'b1010000010100110000010101010000010100000000000001010110000000000,
64'b1100110011000110000000000110110000000110101010101010110000000000,
64'b1010011001100110101010100110000010101100011001101010000011000000,
64'b1010110011000000110001100000000011000110000000001010110011000000,
64'b0000110001100110110011000110000000000110011010100000011000000000,
64'b1100011011000000101010100110000000001100101001100110110001100000,
64'b1010000001101010110000000000000001101100011011001100110011000000,
64'b1010101010100110011001101100000011001010101010101010101001100000,
64'b0110011011001100000000001010000010100110011001100000011010100000,
64'b1010011001101100000010100000000000000000000001101010110011001100,
64'b0110110011001010000000001100000010100110011010101100011000000000,
64'b1010101011001010101001100000000000001100011011000000011001100000,
64'b1010011001101100000010101100000000000000101010100000011000000000,
64'b0110101000001010011001101100000011001100011001100110000011000000,
64'b1100000000000110011001101100000000000000110011001010000010100000,
64'b0110011010101100000010100000000010101100011000001100011011000000,
64'b0000110010101010011011001010000010101100011011000000101001100000,
64'b0000000011001010101000000110000000001100000000000110101010100000,
64'b1100101000000110000010101010101001100110101011000000110011000000,
64'b0110011011000110000001101100000010101010110001101100101011000000,
64'b0000011001101100110000000110000010101010110011000110110000000000,
64'b0110000000000110011010101010000001101100110000001100011000000000,
64'b1100000010101010110010100110000001100000000011000110000001100000,
64'b0110011010100000000000000000000000001100101010100000101001100000,
64'b1010000011001010011011000110000000000000000011001100101001100000,
64'b0000011001100110011011000110000001101010101010101010101001100000,
64'b1100011000001100000010100110000011000000011011000000110011001010,
64'b0110011010100000000001101100000000001010011011000110110010100000,
64'b1010011011001010101011000110000001100000110011001010110011000000,
64'b1100101001101010000000000110000010100000011001101100000000000000,
64'b1010000010100000000001100000000010101010101010100110000001100000,
64'b1010110000001100101011000000000011000000011010100000110000000000,
64'b0110011010100000101000000000000011001010011000001010011001100000,
64'b0000101011000000110010100110000000001010101010101100110001100000,
64'b1010000011001100110010101010110011000110110000001010000000000000,
64'b1100000001101010000001100110000001100110000001100000011010100000,
64'b1010101001101010011000001100000011001100101010100110000010100000,
64'b1010110000001010011000001010000011000000101010101010011000000000,
64'b0000101000000000011001100000000001101010101000000110101011000000,
64'b1100011000001100110011001010000010100000110001101010110001100000,
64'b0000011011001100000001101100000000001010000000000000110001100000,
64'b0110110001100000000010100000000011001100110001100110110001100000,
64'b0000101000000000101011000000000010100000110000000000000010101100,
64'b0110011011000110110001101100000010101100011010101100101001100000,
64'b0000110010100110011000000000000011000000101010100110101000000000,
64'b0000000000001010011011001010000011000000110001100000101010100000,
64'b0110000011001100011011000000000011001100011001100110000011000000,
64'b0000000011000110110000001010000000000000110011001010000010100000,
64'b0000101010101100101010101100000010101100011000001100011011000000,
64'b1010011011001100101011000110000010101100011011000000101001100000,
64'b0110110011000000011010101010000000001100000000000110101010100000,
64'b1010110000001010101001101010101001100110101011000000110011000000,
64'b0110000001101100101000000000000010101010110001101100101011000000,
64'b1010011000000000011011001010000010101010110011000110110000000000,
64'b1010110011000110101001101100000001101100110000001100011000000000,
64'b1010011011001100110001101100000001100000000011000110000001100000,
64'b1100101011001010011000000000000000001100101010100000101001100000,
64'b1010101001100110011001101100000000000000000011001100101001100000,
64'b1010101000001010110010100110000001101010101010101010101001100000,
64'b1100110000000000110011000110000011000000011011000000110011001010,
64'b1100000011001100110000001100000000001010011011000110110010100000,
64'b1010101000001100110010101100000000000000000001101010110011000000,
64'b1100000000000000011010100000000010100000011001101100000000000000,
64'b1010000010100110101010101100000010101010101010100110000001100000,
64'b0000110001101010011011000000000011000000011010100000110000000000,
64'b1100110000001010110000000110000011001010011000001010011001100000,
64'b1100101010101010110001100110000000001010101010101100110001100000,
64'b0110101010101100011011001100110011000110110000001010000000000000,
64'b1100101011000000110010100000000001100110000001100000011010100000,
64'b0110110010101010110000001100000011001100101010100110000010100000,
64'b1100101000001100011001100000000011000000101010101010011000000000,
64'b1100011010101010000001101010000001101010101000000110101011000000,
64'b0000011010100110011010101010000010100000110001101010110001100000,
64'b0110110001101100011011000000000000001010000000000000110001100000,
64'b1100110010100110101001100110000011001100110001100110110001100000,
64'b0000000000000000101000000110000010100000110000000000000010101100,
64'b1010101000000000101010101010000010101100011010101100101001100000,
64'b1100011010100000000011001010000000000000101011000110000010100000,
64'b0000000000001010011011001010000011000000110001100000101010100000,
64'b0110000011001100011011000000000011001100011001100110000011000000,
64'b0000000011000110110000001010000000000000110011001010000010100000,
64'b0000101010101100101010101100000010101100011000001100011011000000,
64'b1010011011001100101011000110000010101100011011000000101001100000,
64'b0110110011000000011010101010000000001100000000000110101010100000,
64'b1010110000001010101001101010101001100110101011000000110011000000,
64'b0110000001101100101000000000000010101010110001101100101011000000,
64'b1010011000000000011011001010000010101010110011000110110000000000,
64'b1010110011000110101001101100000001101100110000001100011000000000,
64'b1010011011001100110001101100000001100000000011000110000001100000,
64'b1100101011001010011000000000000000001100101010100000101001100000,
64'b1010101001100110011001101100000000000000000011001100101001100000,
64'b1010101000001010110010100110000001101010101010101010101001100000,
64'b1100110000000000110011000110000011000000011011000000110011001010,
64'b0000110001101010000010100110000000001010011010100110101001100000,
64'b1010101000001100110010101100000000000000000001101010110011000000,
64'b1100000000000000011010100000000010100000011001101100000000000000,
64'b1010000010100110101010101100000010101010101010100110000001100000,
64'b0000110001101010011011000000000011000000011010100000110000000000,
64'b1100110000001010110000000110000011001010011000001010011001100000,
64'b1100101010101010110001100110000000001010101010101100110001100000,
64'b0110101010101100011011001100110011000110110000001010000000000000,
64'b1100101011000000110010100000000001100110000001100000011010100000,
64'b0110110010101010110000001100000011001100101010100110000010100000,
64'b1100101000001100011001100000000011000000101010101010011000000000,
64'b1100011010101010000001101010000001101010101000000110101011000000,
64'b0000011010100110011010101010000010100000110001101010110001100000,
64'b0110110001101100011011000000000000001010000000000000110001100000,
64'b1100110010100110101001100110000011001100110001100110110001100000,
64'b0000000000000000101000000110000010100000110000000000000010101100,
64'b1010110001101100110010101100101000000110101010101010000010100000,
64'b1100110001101010000000001100000000001100011001100000101010100000,
64'b0110000001101100000001101100000000001010101011001100101000000000,
64'b1010000001100000101011001100000000001100000010101100110000000000,
64'b1100011011001100101011001010000001101010101010100000101000000000,
64'b1100011010100000000011000000000011000110011000001010101000000000,
64'b0000011011000000011011000000000010101010110011001010000000000000,
64'b0000011000001010110011000000000011000000101011001100000000000000,
64'b0110110011001010110010100000000010101010101000001010000000001010,
64'b0110101000000000110000000000000001100110000010101010000000000000,
64'b0110110000000110110000000000000010101100110010100000000000000000,
64'b0110000010101100110000000000000000001010110011000000000000000000,
64'b1100110010101100101000000000000010101010000010100000000010100000,
64'b1010000000001100000000000000000001100000101010100000000000000000,
64'b1100000001101100000000000000000011001100101000000000000000000000,
64'b0000101011001100000000000000000010101100110000000000000000000000,
64'b1100110010100110110001100110110010101100011011001100101001100000,
64'b1100011000001100101000000110000000001010110011000000110011000000,
64'b0000101000001100000010100110000000000110011010100000110000000000,
64'b1100000000001010011001100110000000000000000001101010000000000000,
64'b1100101001101100011001101100000011000110110011001010011000000000,
64'b0110000011001010000001100000000010101100110000001100110000000000,
64'b1010000011000000101001100000000001100110101000001100000000000000,
64'b0000000010100110011001100000000000000000011010100000000000000000,
64'b1010011011000110011011000000000001101100110010100110000000001100,
64'b0000110010100000011000000000000011001100000011001100000000000000,
64'b0000110000001010011000000000000001101010000011000000000000000000,
64'b0000101001100110011000000000000000000110101000000000000000000000,
64'b0110110001100110110000000000000011001100101001100000000011000000,
64'b1100101000000110000000000000000011000000110011000000000000000000,
64'b1100000010100110000000000000000010100000110000000000000000000000,
64'b1010011001100110000000000000000001101010000000000000000000000000,
64'b0000011010100000110011001010000011000000110000001010110011000000,
64'b0110101001100000011010101010101000000110101010101010000010100000,
64'b1100011001100110000010101010000000001100011001100000101010100000,
64'b1010000001100110011000001010000000001010101011001100101000000000,
64'b0110101000001100110010100000000000001100000010101100110000000000,
64'b1010011000000110101010101010000001101010101010100000101000000000,
64'b0110011001100000101010100000000011000110011000001010101000000000,
64'b0000011001100110000010100000000010101010110011001010000000000000,
64'b1010000011001100101000000000000011000000101011001100000000000000,
64'b0110000001101010101010100000000010101010101000001010000000001010,
64'b0110011000001010101000000000000001100110000010101010000000000000,
64'b0110011001100000101000000000000010101100110010100000000000000000,
64'b0000110011001010000000000000000000001010110011000000000000000000,
64'b0000011010101010101000000000000010101010000010100000000010100000,
64'b0110000010101010000000000000000001100000101010100000000000000000,
64'b0110011000001010000000000000000011001100101000000000000000000000,
64'b1010110011001010101010101100000000000000000000000110101000000000,
64'b1100011011000000011001101100110010101100011011001100101001100000,
64'b1010110001101100101011001100000000001010110011000000110011000000,
64'b0110101001100110110000001100000000000110011010100000110000000000,
64'b1100110010101010101011000000000000000000000001101010000000000000,
64'b0110110000000110011011001100000011000110110011001010011000000000,
64'b1100011011001010110011000000000010101100110000001100110000000000,
64'b1010011001101100000011000000000001100110101000001100000000000000,
64'b1100101010101010110000000000000000000000011010100000000000000000,
64'b1100000001100110110011000000000001101100110010100110000000001100,
64'b0110110010101100110000000000000011001100000011001100000000000000,
64'b0110011011000000110000000000000001101010000011000000000000000000,
64'b1010101010101100000000000000000000000110101000000000000000000000,
64'b0000011001101100110000000000000011001100101001100000000011000000,
64'b1100101011001100000000000000000011000000110011000000000000000000,
64'b0110110000001100000000000000000010100000110000000000000000000000,
64'b1100011001101010101011001100000000000000101010101100110010100000,
64'b1100101011001010110011000110000011000000110000001010110011000000,
64'b0000101000001100011011000110101000000110101010101010000010100000,
64'b0110011000000110101001100110000000001100011001100000101010100000,
64'b0110011010101010110011000000000000001010101011001100101000000000,
64'b1010110010101100110001100000000000001100000010101100110000000000,
64'b1010000011000110110001101010000001101010101010100000101000000000,
64'b0110000001101010011001100000000011000110011000001010101000000000,
64'b0110101010101100110000000000000010101010110011001010000000000000,
64'b1100101011001100011000000000000011000000101011001100000000000000,
64'b0000110001101100011010100000000010101010101000001010000000001010,
64'b0000011010100110011000000000000001100110000010101010000000000000,
64'b1010101011001100000000000000000010101100110010100000000000000000,
64'b1010110011000110000000000000000000001010110011000000000000000000,
64'b1100011011000110101000000000000010101010000010100000000010100000,
64'b0110101001100110000000000000000001100000101010100000000000000000,
64'b1010101000000000101010100110000000000000011001101010000011000000,
64'b0110101011000110000010101010000000000000000000000110101000000000,
64'b1100110011001100011011001010110010101100011011001100101001100000,
64'b0110110001100110110010101010000000001010110011000000110011000000,
64'b1010000000001010101001100000000000000110011010100000110000000000,
64'b1010110001100000101010100000000000000000000001101010000000000000,
64'b1100110011000110110010101100000011000110110011001010011000000000,
64'b1100011001101100101010100000000010101100110000001100110000000000,
64'b0000000010101010011000000000000001100110101000001100000000000000,
64'b1100011000001010101000000000000000000000011010100000000000000000,
64'b1100110001101100101011000000000001101100110010100110000000001100,
64'b0110011011001010101000000000000011001100000011001100000000000000,
64'b0000101010100110000000000000000001101010000011000000000000000000,
64'b0110000010101010000000000000000000000110101000000000000000000000,
64'b1100011011001010110000000000000011001100101001100000000011000000,
64'b0110110010101010000000000000000011000000110011000000000000000000,
64'b0110011010101010011001101100000010101100101010101010101001100000,
64'b1100110000001100000011000110000011001100110000001100110001100000,
64'b1010000010101010110000001100000010100000101011001010101000000000,
64'b0110101001100110101001101100101010100110110010100000110001100000,
64'b0110101010100110011011000000000011001010101010101010011000000000,
64'b1100000011000000110001100000000011001100000011001100011000000000,
64'b0000101010101100000011000000000000001010110010101010000000000000,
64'b1010011001101010011011001010000001101100101000001100011000000000,
64'b1010101001100110110000000000000010101010101010100110000000000000,
64'b0000110000001100011000000000000011000000110011000110000000000000,
64'b1010101011000000110000000000000010101100101010100000000000000000,
64'b0110011010100110110010100000000011001010000011000110000000001010,
64'b1010011001101100000000000000000010101010101001100000000000000000,
64'b1100000011000110000000000000000000001100110001100000000000000000,
64'b1010110000001100000000000000000011001010101000000000000000000000,
64'b0110101001101100101000000000000010100000110001100000000010100000,
64'b0110101010101010101001100110000011001100000010100000011010100000,
64'b0110011001101010101010101010000011000110011010100000000010100000,
64'b0000101010101010000011000110000000001010000011000110000001100000,
64'b0110110010101100110000000110110001101100011001101010110000000000,
64'b1010101010101010011001100000000011000000101000000110101000000000,
64'b0110011010101010101010100000000001100110101000000000101000000000,
64'b1010101010100000110001100000000010100000110001100000011000000000,
64'b1100101011001100000001101100000011000110011010101100000000000000,
64'b1010101010100110011000000000000000001010000001101010000000000000,
64'b0110101010101010101000000000000001101010000000001010000000000000,
64'b1010101000001100011000000000000000001100011000000110000000000000,
64'b1010110011000000011011000000000001100110101011000000000000001100,
64'b1010101001100110000000000000000010100000011010100000000000000000,
64'b1010101010101010000000000000000010100000000010100000000000000000,
64'b1010000011000110000000000000000011000110000001100000000000000000,
64'b1100110000000110110000000000000001101010110000000000000011000000,
64'b0110101000000000101011000000000000001010101001101010110001100000,
64'b1010000010100110110001101010000010100110110011000000101011000000,
64'b1100011000000000000001100000000010100110101000001100000011000000,
64'b0110000010100000101001101010000011000000110001100110000010100000,
64'b1010000000001010110000000000101010101010011010101100011000000000,
64'b0000101001101100011010100000000001101100110000001010110000000000,
64'b0110000000000000011000000000000001101010000011000000110000000000,
64'b0000101000001010011010100000000000001100011001100000101000000000,
64'b0000000010101100000000001010000010100110101011000110000000000000,
64'b1010011011000110101000000000000011001100000010101100000000000000,
64'b0000000000000110000000000000000010100000110000001100000000000000,
64'b1010000010100110101000000000000011000110011000001010000000000000,
64'b0000101011000000000010100000000001101010110001100000000000001010,
64'b0110110001101010000000000000000011000000101011000000000000000000,
64'b0000000001100000000000000000000000001100000011000000000000000000,
64'b0000101001101010000000000000000001100110000010100000000000000000,
64'b0110011000000000110000001010000000000110110001100110101011000000,
64'b0110000011001100000001101100000011001100000010100000011010100000,
64'b0000110000001010101001100000000011000110011010100000000010100000,
64'b0110101011000000110001101100000000001010000011000110000001100000,
64'b0110000000001100000010100000110001101100011001101010110000000000,
64'b0000110011000000011011000000000011000000101000000110101000000000,
64'b1100000010101010011000000000000001100110101000000000101000000000,
64'b1010110000001100011011000000000010100000110001100000011000000000,
64'b0000000011000000101000001100000011000110011010101100000000000000,
64'b1100110000000110110000000000000000001010000001101010000000000000,
64'b0000101010100110000000000000000001101010000000001010000000000000,
64'b1100000011000110110000000000000000001100011000000110000000000000,
64'b0000110000001010000011000000000001100110101011000000000000001100,
64'b1100000001101100000000000000000010100000011010100000000000000000,
64'b1010101001100000000000000000000010100000000010100000000000000000,
64'b0000110001101100000000000000000011000110000001100000000000000000,
64'b0110101001100110110000001010000010100000011000001010110011000000,
64'b1010011001101010101011001100000011000110110011001010110010100000,
64'b1100000011001010110000000110000011000110101000000000110000000000,
64'b0110011001100000101010101100000000000110110000000110110000000000,
64'b1010011001101100000010100000000000000110000010101100110000000000,
64'b0110011010101010110011000000101001101100110010101100101000000000,
64'b0000110010101100000001100000000001101010000000001100000000000000,
64'b0110011000001010101011000000000001101100000001101100000000000000,
64'b0110011011000000101000000000000001100000101011001100000000000000,
64'b0110101010101100110000001010000011001100101011001010000000000000,
64'b1100101011000000011000000000000010100000000011000000000000000000,
64'b0110000010101010110000000000000011000000011011000000000000000000,
64'b0110110000001010000000000000000000001010110011000000000000000000,
64'b1010101011001100000010100000000011001010110010100000000000001010,
64'b1010110000000110000000000000000000000000110000000000000000000000,
64'b0000101010101100000000000000000000000110110000000000000000000000,
64'b0110101000001010110010100000000001100000011010101100101010100000,
64'b1010000000001100011000001100000000001100101000001100101001100000,
64'b0110101011000000000011001010000010100110011010100000101000000000,
64'b1100110000000000110000000110000010100110000000001100101000000000,
64'b1010000010101100101000000000000000000110101011001010101000000000,
64'b0000000011000110000011000000110011001010000011001010011000000000,
64'b1010110000000000110010100000000001100110101000001010000000000000,
64'b1100000000001100000001100000000001100000000011001010000000000000,
64'b0000101011001010000000000000000001101010110010101010000000000000,
64'b0000110001100000110000001100000010100000110010100110000000000000,
64'b1100000000001100101000000000000001101010000010100000000000000000,
64'b0000000011000000011000000000000000000000110010100000000000000000,
64'b1010110010100000000000000000000010101100101010100000000000000000,
64'b1100011000001100000011000000000000001100101001100000000000001100,
64'b0000000011001010000000000000000010100000101000000000000000000000,
64'b0000110000000110000000000000000000001100101000000000000000000000,
64'b0110101011000000110011001100000001100000011011000000011011000000,
64'b1010110001101010011000001100000010100000011000001010110011000000,
64'b1010110001100110101001101010000011000110110011001010110010100000,
64'b0000000011000000101001100000000011000110101000000000110000000000,
64'b1010110000001100110011000000000000000110110000000110110000000000,
64'b1100011010100110000011000000000000000110000010101100110000000000,
64'b1100011001101010011010100000101001101100110010101100101000000000,
64'b0000110000001010011000000000000001101010000000001100000000000000,
64'b1100000011001100110000000000000001101100000001101100000000000000,
64'b0110101001100000110000000000000001100000101011001100000000000000,
64'b0110011010100110101000001010000011001100101011001010000000000000,
64'b1100000010100110000000000000000010100000000011000000000000000000,
64'b0000110011001100000000000000000011000000011011000000000000000000,
64'b1010011000001100000000000000000000001010110011000000000000000000,
64'b0110101001101010000010100000000011001010110010100000000000001010,
64'b0000101001100000000000000000000000000000110000000000000000000000,
64'b0110110000001010000000001010000001101010011000000000110010100000,
64'b0110000001101100011010101010000001100000011010101100101010100000,
64'b1100101001101100011011000110000000001100101000001100101001100000,
64'b0000101010101010110001100000000010100110011010100000101000000000,
64'b1100000010100000000010100000000010100110000000001100101000000000,
64'b0000011011000110101010100000000000000110101011001010101000000000,
64'b1010011011000110110001100000110011001010000011001010011000000000,
64'b1010101010101100011000000000000001100110101000001010000000000000,
64'b0000101000000000101000000000000001100000000011001010000000000000,
64'b0110110001101010101000000000000001101010110010101010000000000000,
64'b0110110001101100011000001100000010100000110010100110000000000000,
64'b1010101011000110000000000000000001101010000010100000000000000000,
64'b1010000000001010000000000000000000000000110010100000000000000000,
64'b1100011010101010000000000000000010101100101010100000000000000000,
64'b1100011011000110000011000000000000001100101001100000000000001100,
64'b1010110001100000000000000000000010100000101000000000000000000000,
64'b1100000000001100000010100110000011001100011010100000000011000000,
64'b0110101011000000110011001100000001100000011011000000011011000000,
64'b1010110001101010011000001100000010100000011000001010110011000000,
64'b1010110001100110101001101010000011000110110011001010110010100000,
64'b0000000011000000101001100000000011000110101000000000110000000000,
64'b1010110000001100110011000000000000000110110000000110110000000000,
64'b1100011010100110000011000000000000000110000010101100110000000000,
64'b1100011001101010011010100000101001101100110010101100101000000000,
64'b0000110000001010011000000000000001101010000000001100000000000000,
64'b1100000011001100110000000000000001101100000001101100000000000000,
64'b0110101001100000110000000000000001100000101011001100000000000000,
64'b0110011010100110101000001010000011001100101011001010000000000000,
64'b1100000010100110000000000000000010100000000011000000000000000000,
64'b0000110011001100000000000000000011000000011011000000000000000000,
64'b1010011000001100000000000000000000001010110011000000000000000000,
64'b0110101001101010000010100000000011001010110010100000000000001010,
64'b0000000010101010101011000110000000001010011001101010000010100000,
64'b0110110000001010000000001010000001101010011000000000110010100000,
64'b0110000001101100011010101010000001100000011010101100101010100000,
64'b1100101001101100011011000110000000001100101000001100101001100000,
64'b0000101010101010110001100000000010100110011010100000101000000000,
64'b1100000010100000000010100000000010100110000000001100101000000000,
64'b0000011011000110101010100000000000000110101011001010101000000000,
64'b1010011011000110110001100000110011001010000011001010011000000000,
64'b1010101010101100011000000000000001100110101000001010000000000000,
64'b0000101000000000101000000000000001100000000011001010000000000000,
64'b0110110001101010101000000000000001101010110010101010000000000000,
64'b0110110001101100011000001100000010100000110010100110000000000000,
64'b1010101011000110000000000000000001101010000010100000000000000000,
64'b1010000000001010000000000000000000000000110010100000000000000000,
64'b1100011010101010000000000000000010101100101010100000000000000000,
64'b1100011011000110000011000000000000001100101001100000000000001100

};

parameter [0:12287] C_POLY =  
{
64'h55555555aaaaaaaa,
64'h6699669999669966,
64'h6699996666999966,
64'h9966669966999966,
64'hcc3333cccc3333cc,
64'hf0f0f0f0f0f0f0f0,
64'h33333333cccccccc,
64'h0ff0f00ff00f0ff0,
64'hf00ff00f0ff00ff0,
64'ha55aa55aa55aa55a,
64'h9669966969966996,
64'hf0f0f0f0f0f0f0f0,
64'h0f0f0f0ff0f0f0f0,
64'h3333cccc3333cccc,
64'hcccccccccccccccc,
64'hffffffff00000000,
64'hf0f0f0f0f0f0f0f0,
64'h5a5a5a5a5a5a5a5a,
64'hff00ff00ff00ff00,
64'ha5a5a5a55a5a5a5a,
64'hf0f0f0f0f0f0f0f0,
64'h0000000000000000,
64'h55aa55aa55aa55aa,
64'h3c3c3c3c3c3c3c3c,
64'haaaa55555555aaaa,
64'h55555555aaaaaaaa,
64'h3333cccc3333cccc,
64'h9966669966999966,
64'hff00ff00ff00ff00,
64'hf0f0f0f0f0f0f0f0,
64'h6666666666666666,
64'h00ff00ffff00ff00,
64'hc33c3cc33cc3c33c,
64'ha55aa55aa55aa55a,
64'h9966996699669966,
64'hf0f0f0f0f0f0f0f0,
64'h9696969696969696,
64'hffff0000ffff0000,
64'ha55a5aa55aa5a55a,
64'h6699996666999966,
64'hc3c33c3cc3c33c3c,
64'hf0f0f0f0f0f0f0f0,
64'h3cc33cc3c33cc33c,
64'h9966996699669966,
64'h55555555aaaaaaaa,
64'h0ff00ff00ff00ff0,
64'h3c3cc3c3c3c33c3c,
64'hf0f0f0f0f0f0f0f0,
64'h0ff0f00ff00f0ff0,
64'h0ff0f00ff00f0ff0,
64'haa5555aaaa5555aa,
64'h33333333cccccccc,
64'h3c3cc3c3c3c33c3c,
64'h5a5a5a5a5a5a5a5a,
64'h55aaaa55aa5555aa,
64'h55aaaa55aa5555aa,
64'h6666999999996666,
64'hf0f0f0f0f0f0f0f0,
64'h5aa55aa5a55aa55a,
64'h9696969696969696,
64'h9999666699996666,
64'h00ffff0000ffff00,
64'h0ff0f00ff00f0ff0,
64'hcccc33333333cccc,
64'h0000000000000000,
64'h9696969696969696,
64'h9696969696969696,
64'h6699996666999966,
64'h9999999966666666,
64'h3cc3c33c3cc3c33c,
64'h6699996666999966,
64'h3c3c3c3c3c3c3c3c,
64'h9669966969966996,
64'h5aa5a55a5aa5a55a,
64'h5aa5a55a5aa5a55a,
64'h3c3c3c3c3c3c3c3c,
64'hf00ff00f0ff00ff0,
64'hf0f0f0f0f0f0f0f0,
64'h9669699696696996,
64'h9966669966999966,
64'h33cccc33cc3333cc,
64'h0ff00ff00ff00ff0,
64'h00ffff0000ffff00,
64'h5a5a5a5a5a5a5a5a,
64'h6996966996696996,
64'h3c3cc3c3c3c33c3c,
64'h5a5aa5a5a5a55a5a,
64'haa5555aaaa5555aa,
64'h0000ffffffff0000,
64'h3c3c3c3c3c3c3c3c,
64'hc33c3cc33cc3c33c,
64'h5aa55aa5a55aa55a,
64'h6699669999669966,
64'h6666999999996666,
64'hffffffff00000000,
64'h5a5a5a5a5a5a5a5a,
64'h5aa5a55a5aa5a55a,
64'h0000ffffffff0000,
64'h0ff00ff00ff00ff0,
64'hf00f0ff0f00f0ff0,
64'h6699996666999966,
64'h9696969696969696,
64'h33cccc33cc3333cc,
64'hffffffff00000000,
64'haa5555aaaa5555aa,
64'hff0000ff00ffff00,
64'h3c3cc3c3c3c33c3c,
64'h3c3c3c3c3c3c3c3c,
64'h5a5aa5a5a5a55a5a,
64'haaaaaaaaaaaaaaaa,
64'h6666999999996666,
64'h0000ffffffff0000,
64'h5aa55aa5a55aa55a,
64'h5a5a5a5a5a5a5a5a,
64'hcc33cc3333cc33cc,
64'h6666666666666666,
64'hc3c3c3c33c3c3c3c,
64'h55555555aaaaaaaa,
64'h6699996666999966,
64'h9696969696969696,
64'h0f0ff0f00f0ff0f0,
64'h9696969696969696,
64'h0ff00ff00ff00ff0,
64'h6666666666666666,
64'h9696696969699696,
64'h3c3c3c3c3c3c3c3c,
64'h00ff00ffff00ff00,
64'hc33cc33cc33cc33c,
64'h00ffff0000ffff00,
64'h3c3c3c3c3c3c3c3c,
64'h3cc33cc3c33cc33c,
64'h5a5a5a5a5a5a5a5a,
64'h0000ffffffff0000,
64'h3c3cc3c3c3c33c3c,
64'h6699669999669966,
64'h9696696969699696,
64'h3c3c3c3c3c3c3c3c,
64'h9696969696969696,
64'haaaaaaaaaaaaaaaa,
64'h3c3c3c3c3c3c3c3c,
64'h0ff00ff00ff00ff0,
64'h0f0ff0f00f0ff0f0,
64'h6969969669699696,
64'h3c3c3c3c3c3c3c3c,
64'hcccccccccccccccc,
64'h0ff00ff00ff00ff0,
64'h00ffff0000ffff00,
64'h00ff00ffff00ff00,
64'h3cc33cc3c33cc33c,
64'hf0f0f0f0f0f0f0f0,
64'h5a5a5a5a5a5a5a5a,
64'h00ffff0000ffff00,
64'h0000ffffffff0000,
64'hffff0000ffff0000,
64'h5aa5a55a5aa5a55a,
64'h5a5a5a5a5a5a5a5a,
64'h6699669999669966,
64'h6699996666999966,
64'h9966669966999966,
64'hcc3333cccc3333cc,
64'hffffffff00000000,
64'h3c3c3c3c3c3c3c3c,
64'h6969969669699696,
64'h9696696969699696,
64'h3c3cc3c3c3c33c3c,
64'h5a5aa5a5a5a55a5a,
64'h0000000000000000,
64'h5a5a5a5a5a5a5a5a,
64'h3cc33cc3c33cc33c,
64'h3cc33cc3c33cc33c,
64'h5aa55aa5a55aa55a,
64'h6699669999669966,
64'haaaaaaaaaaaaaaaa,
64'h3c3c3c3c3c3c3c3c,
64'hf00f0ff0f00f0ff0,
64'h5aa5a55a5aa5a55a,
64'h6699996666999966,
64'h6969969669699696,
64'h6666666666666666,
64'hf0f0f0f0f0f0f0f0,
64'hff0000ff00ffff00,
64'h33cccc33cc3333cc,
64'h3c3cc3c3c3c33c3c,
64'h3cc33cc3c33cc33c,
64'h3c3c3c3c3c3c3c3c,
64'hf0f0f0f0f0f0f0f0,
64'h0000ffffffff0000,
64'h5a5aa5a5a5a55a5a,
64'h5aa55aa5a55aa55a,
64'h5aa5a55a5aa5a55a,
64'ha55aa55aa55aa55a,
64'hf0f0f0f0f0f0f0f0
};

parameter [1023:0] AHEAD_POLY = { 
32'b10000111010111011011011101011000,
32'b01000100111100110110110011110100,
32'b00100101001001000000000100100010,
32'b00010010100100100000000010010001,
32'b10001110000101001011011100010000,
32'b11000000010101111110110011010000,
32'b11100000001010111111011001101000,
32'b01110111010010000100110001101100,
32'b00111100111110011001000101101110,
32'b10011110011111001100100010110111,
32'b11001000011000111101001100000011,
32'b11100011011011000101111011011001,
32'b11110110111010111001100000110100,
32'b11111011011101011100110000011010,
32'b11111101101110101110011000001101,
32'b01111110110111010111001100000110,
32'b10111000001100110000111011011011,
32'b01011100000110011000011101101101,
32'b10101110000011001100001110110110,
32'b01010111000001100110000111011011,
32'b00101011100000110011000011101101,
32'b00010101110000011001100001110110,
32'b00001101101111010111101101100011,
32'b10000001100000110000101011101001,
32'b01000000110000011000010101110100,
32'b10100000011000001100001010111010,
32'b11010111011011011101011000000101,
32'b11101011101101101110101100000010,
32'b01110101110110110111010110000001,
32'b00111010111011011011101011000000,
32'b00011101011101101101110101100000,
32'b00001110101110110110111010110000

  } ;




//*******************
//DEFINE LOCAL PARAMETER
//*******************
//parameter(s)

 wire              crc_en_pre ;
 wire  [31:0]      crc_pre    ;

function [7:0] reverse_8b;
  input [7:0]   data;
  integer        k;
    begin
        for (k = 0; k < 8; k = k + 1) begin
            reverse_8b[k] = data[7 - k];
        end
    end
endfunction

// 定义对数函数  来自https://blog.csdn.net/w40306030072/article/details/79014822，并修改
function integer clogb2 (input integer bit_depth);
begin
for(clogb2=0; bit_depth>1; clogb2=clogb2+1)
bit_depth = bit_depth>>1;
end
endfunction
 

//*********************
//INNER SIGNAL DECLARATION
//*********************
//REGS
  

//WIRES
// wire [31:0] crc_pipe;

// wire                 sop_lut_pipe  ;
// wire                 eop_lut_pipe  ;
// wire                dval_lut_pipe  ;
// wire [MOD_WIDTH:0]   mod_lut_pipe  ;
// wire [31:0]         dout_lut_pipe  ;

wire  [SEG_NUM-1:0]            lut_pipe_sop_out        ;
wire  [SEG_NUM-1:0]            lut_pipe_eop_out        ;
wire  [SEG_NUM-1:0]            lut_pipe_dval_out       ;
wire  [SEG_NUM*4-1:0]          lut_pipe_packet_num_out ;
wire  [SEG_NUM*12-1:0]         lut_pipe_zero_num_out   ;
wire  [SEG_NUM*32-1:0]         lut_pipe_dout_out       ;



//*********************
//INSTANTCE MODULE
//*********************

// lut_pipe_top  u_lut_pipe_top   (     
//         .clk       ( clk      )   ,
//         .rst       ( rst      )   ,
//         .din_en    ( dval     )   ,
//         .din       ( din      )   ,
//         .dout      ( crc_pipe )    
//               ) ;

// wire [31:0] crc_pipe_new ;

  lut_pipe_multi   

# ( 

    .D_LUT_POLY            ( D_LUT_POLY          ) ,
    .D_CRC_REG_INIT        ( D_CRC_REG_INIT        ) ,
    .SEG_NUM             ( SEG_NUM             )  ,
    .BUS_WIDTH           ( BUS_WIDTH           )  ,
    .BUS_WIDTH_MULTI_6   ( BUS_WIDTH_MULTI_6   )  ,
    .MOD_WIDTH           ( MOD_WIDTH           )  ,
    .CMP_LAYER           ( CMP_LAYER           )  ,      // C_XOR之前计算的层数，包含第一层
    .LUT_NUM_LAYER_1     ( LUT_NUM_LAYER_1     )  ,
    .LUT_NUM_LAYER_2     ( LUT_NUM_LAYER_2     )  ,
    .LUT_NUM_LAYER_3     ( LUT_NUM_LAYER_3     )  ,
    .LUT_NUM_LAYER_4     ( LUT_NUM_LAYER_4     )  ,
    .LUT_NUM_LAYER_5     ( LUT_NUM_LAYER_5     )  ,
    .LUT_NUM_LAYER_6     ( LUT_NUM_LAYER_6     )  ,
    .LUT_NUM_LAYER_7     ( LUT_NUM_LAYER_7     )  ,
    .LUT_NUM_LAYER_8     ( LUT_NUM_LAYER_8     )  ,        
    .LUT_OUT_NUM_LAYER_1 ( LUT_OUT_NUM_LAYER_1 )  ,
    .LUT_OUT_NUM_LAYER_2 ( LUT_OUT_NUM_LAYER_2 )  ,
    .LUT_OUT_NUM_LAYER_3 ( LUT_OUT_NUM_LAYER_3 )  ,
    .LUT_OUT_NUM_LAYER_4 ( LUT_OUT_NUM_LAYER_4 )  ,
    .LUT_OUT_NUM_LAYER_5 ( LUT_OUT_NUM_LAYER_5 )  ,
    .LUT_OUT_NUM_LAYER_6 ( LUT_OUT_NUM_LAYER_6 )  ,
    .LUT_OUT_NUM_LAYER_7 ( LUT_OUT_NUM_LAYER_7 )  ,
    .LUT_OUT_NUM_LAYER_8 ( LUT_OUT_NUM_LAYER_8 )      

  ) u_lut_pipe_multi
(     
    .clk       ( clk     ) ,
    .rst       ( rst     ) ,

    .seg_sop        ( seg_sop        ) ,
    .seg_eop        ( seg_eop        ) ,
    .seg_dval       ( seg_dval       ) ,
    .seg_packet_num ( seg_packet_num ) ,
    .seg_zero_num   ( seg_zero_num   ) ,
    .seg_dout       ( seg_dout       ) ,

    

    .sop_out        ( lut_pipe_sop_out        )  ,
    .eop_out        ( lut_pipe_eop_out        )  ,
    .dval_out       ( lut_pipe_dval_out       )  ,
    .packet_num_out ( lut_pipe_packet_num_out )  ,
    .zero_num_out   ( lut_pipe_zero_num_out   )  ,
    .dout_out       ( lut_pipe_dout_out       )   

              ) ;



wire  [PKT_NUM-1:0]           merge_eop_out        ;
wire  [PKT_NUM-1:0]           merge_dval_out       ;
wire  [4 *( PKT_NUM )-1:0]    merge_packet_num_out ;
wire  [12*( PKT_NUM )-1:0]    merge_zero_num_out   ;
wire  [32*( PKT_NUM )-1:0]    merge_dout_out       ;

merge_top 

# ( 
        .SEG_NUM    ( SEG_NUM    ),
        .AHEAD_POLY ( AHEAD_POLY ),
        .PKT_NUM    ( PKT_NUM ) // 1 个最短包512bit 

  ) 

u_merge_top ( 

       . clk ( clk ) ,
       . rst ( rst ) ,
       . lut_pipe_sop_out        ( lut_pipe_sop_out        ) ,        
       . lut_pipe_eop_out        ( lut_pipe_eop_out        ) ,
       . lut_pipe_dval_out       ( lut_pipe_dval_out       ) ,
       . lut_pipe_packet_num_out ( lut_pipe_packet_num_out ) ,
       . lut_pipe_zero_num_out   ( lut_pipe_zero_num_out   ) ,
       . lut_pipe_dout_out       ( lut_pipe_dout_out       ) ,

       .  merge_eop_out         ( merge_eop_out        ) ,
       .  merge_dval_out        ( merge_dval_out       ) ,
       .  merge_packet_num_out  ( merge_packet_num_out ) ,
       .  merge_zero_num_out    ( merge_zero_num_out   ) ,
       .  merge_dout_out        ( merge_dout_out       ) 



 ) ;


// wire  [PKT_NUM-1:0]           t_crossbar_64_merge_sop_out        ;
// wire  [PKT_NUM-1:0]           t_crossbar_64_merge_eop_out        ;
// wire  [PKT_NUM-1:0]           t_crossbar_64_merge_dval_out       ;
// wire  [4 *( PKT_NUM )-1:0]    t_crossbar_64_merge_packet_num_out ;
// wire  [12*( PKT_NUM )-1:0]    t_crossbar_64_merge_zero_num_out   ;
// wire  [32*( PKT_NUM )-1:0]    t_crossbar_64_merge_dout_out       ;

c_xor_and_go_back_top  

 # (              
         .GO_BACK_STAGE ( GO_BACK_STAGE )   ,
         .PKT_NUM       ( PKT_NUM       )   ,
         .GO_BACK_POLY  ( GO_BACK_POLY_STRIDE_8  )   ,
         .C_POLY        ( C_POLY )  
   ) u_c_xor_and_go_back_top
( 
            .clk ( clk )  ,
            .rst ( rst )  ,

            .eop_in  (  merge_eop_out   ) ,  //         // t_crossbar_64_merge_eop_out
            .dval_in (  merge_dval_out   ) ,  //        // t_crossbar_64_merge_dval_out
            .mod_in  (  merge_zero_num_out   ) ,  //    // t_crossbar_64_merge_zero_num_out
            .din     (  merge_dout_out   ) ,  //        // t_crossbar_64_merge_dout_out
                     
            .crc_en_out  ( crc_en ) ,
            .crc_out     ( crc    )


 ) ;







 







//*********************
//MAIN CORE
//********************* 


// always @(posedge clk or posedge rst) begin
//     if (rst) begin
//         crc_en <= 'b0  ;
//         crc    <= 'b0  ;
//     end
//     else begin
//         crc_en <= crc_en_pre  ;
//         crc    <= // crc_pre ;
//                 {  ~reverse_8b(crc_pre[31:24]) ,  
//                    ~reverse_8b(crc_pre[23:16]) ,  
//                    ~reverse_8b(crc_pre[15:8])  , 
//                    ~reverse_8b(crc_pre[7:0])
//                } ; 
//     end
// end

// always @(posedge clk or posedge rst) begin
//     if (rst) begin
//         crc_en <= 'b0  ;
//         crc    <= 'b0  ;
//     end
//     else begin
//         crc_en <= crc_en_pre  ;
//         crc    <=  crc_pre ;
//     end
// end


// always @(posedge clk or posedge rst) begin
//     if (rst) begin
//         crc_en <= 'b0  ;
//         crc    <= 'b0  ;
//     end
//     else begin
//         crc_en <= merge_eop_out  ;
//         crc    <=  merge_dout_out ;
//     end
// end



// test : see merge out ========================================================================


// reg            out_see_merge_eop_out[0:7]   ;
// reg            out_see_merge_dval_out[0:7]  ;
// reg [3:0]      out_see_merge_packet_num_out[0:7] ; // 4bit*64seg
// reg [11:0]     out_see_merge_zero_num_out[0:7] ; // 12bit*64seg the bytes from eo(in a certain segment) to the end of the beat(some segment are treated aszeros); 单位是字节
// reg [31:0]     out_see_merge_dout_out[0:7]  ; // 4096 bits with 64 seg  

// integer k ;
// always @(*) begin

//     for ( k=0; k<8; k=k+1 ) begin
//                out_see_merge_eop_out[k] <=  merge_eop_out [k]                              ;
//               out_see_merge_dval_out[k] <=  merge_dval_out[k]                              ;
//         out_see_merge_packet_num_out[k] <=  merge_packet_num_out [k*4+3 -: 4   ] ;
//           out_see_merge_zero_num_out[k] <=  merge_zero_num_out   [k*12+11 -: 12] ;
//               out_see_merge_dout_out[k] <=  merge_dout_out       [(k+1)*32-1 -: 32] ;
//     end


// end


// test 64*64 crossbar ==================================================================
// wire  [PKT_NUM-1:0]           crossbar_64_merge_sop_out        ;
// wire  [PKT_NUM-1:0]           crossbar_64_merge_eop_out        ;
// wire  [PKT_NUM-1:0]           crossbar_64_merge_dval_out       ;
// wire  [4 *( PKT_NUM )-1:0]    crossbar_64_merge_packet_num_out ;
// wire  [12*( PKT_NUM )-1:0]    crossbar_64_merge_zero_num_out   ;
// wire  [32*( PKT_NUM )-1:0]    crossbar_64_merge_dout_out       ;




// merge_crossbar 

// # ( 

//     .SEG_NUM_IN  ( 64 ) , // 8 in
//     .PKT_NUM_OUT ( 8 )   // 8 out
//   )

// u_merge_crossbar    ( 

//         .clk ( clk ) ,
//         .rst ( rst ) ,

//         .in_sop        ( lut_pipe_sop_out         ) ,
//         .in_eop        ( lut_pipe_eop_out         ) ,
//         .in_dval       ( lut_pipe_dval_out        ) ,
//         .in_packet_num ( lut_pipe_packet_num_out  ) ,
//         .in_zero_num   ( lut_pipe_zero_num_out    ) ,
//         .in_dout       ( lut_pipe_dout_out        ) ,

//         .out_sop        ( crossbar_64_merge_sop_out         ) ,
//         .out_eop        ( crossbar_64_merge_eop_out         ) ,
//         .out_dval       ( crossbar_64_merge_dval_out        ) ,
//         .out_packet_num ( crossbar_64_merge_packet_num_out  ) ,
//         .out_zero_num   ( crossbar_64_merge_zero_num_out    ) ,
//         .out_dout       ( crossbar_64_merge_dout_out        )



//  ) ;


// reg            c_out_see_merge_eop_out[0:7]   ;
// reg            c_out_see_merge_dval_out[0:7]  ;
// reg [3:0]      c_out_see_merge_packet_num_out[0:7] ; // 4bit*64seg
// reg [11:0]     c_out_see_merge_zero_num_out[0:7] ; // 12bit*64seg the bytes from eo(in a certain segment) to the end of the beat(some segment are treated aszeros); 单位是字节
// reg [31:0]     c_out_see_merge_dout_out[0:7]  ; // 4096 bits with 64 seg  

// integer kkk ;
// always @(*) begin

//     for ( kkk=0; kkk<8; kkk=kkk+1 ) begin
//                c_out_see_merge_eop_out[kkk] <=  crossbar_64_merge_eop_out [kkk]                              ;
//               c_out_see_merge_dval_out[kkk] <=  crossbar_64_merge_dval_out[kkk]                              ;
//         c_out_see_merge_packet_num_out[kkk] <=  crossbar_64_merge_packet_num_out [kkk*4+3 -: 4   ] ;
//           c_out_see_merge_zero_num_out[kkk] <=  crossbar_64_merge_zero_num_out   [kkk*12+11 -: 12] ;
//               c_out_see_merge_dout_out[kkk] <=  crossbar_64_merge_dout_out       [(kkk+1)*32-1 -: 32] ;
//     end


// end



// assign t_crossbar_64_merge_eop_out       = crossbar_64_merge_eop_out      ;
// assign t_crossbar_64_merge_dval_out      = crossbar_64_merge_dval_out     ;
// assign t_crossbar_64_merge_zero_num_out  = crossbar_64_merge_zero_num_out ;
// assign t_crossbar_64_merge_dout_out      = crossbar_64_merge_dout_out     ;


// test merge module ==============================================================







// reg              seri_lut_pipe_eop_out         [0:SEG_NUM-1]    ;
// reg              seri_lut_pipe_dval_out        [0:SEG_NUM-1]    ;
// reg  [3:0]       seri_lut_pipe_packet_num_out  [0:SEG_NUM-1]    ;
//        // wire  [11:0]      seri_lut_pipe_zero_num_out    [0:SEG_NUM-1]    ;
// reg  [31:0]      seri_lut_pipe_dout_out        [0:SEG_NUM-1]    ;


// integer ii ;

// always @(*) begin

//     for ( ii=0; ii<64; ii=ii+1 ) begin
//                  seri_lut_pipe_eop_out        [ii]     <=   lut_pipe_eop_out         [ii]                      ;
//                  seri_lut_pipe_dval_out       [ii]     <=   lut_pipe_dval_out        [ii]                      ;
//                  seri_lut_pipe_packet_num_out [ii]     <=   lut_pipe_packet_num_out  [ii*4+3 -: 4   ]          ;
//                  // seri_lut_pipe_zero_num_out   [ii]     <=   lut_pipe_zero_num_out    [ii*12+11 -: 12]          ;
//                  seri_lut_pipe_dout_out       [ii]     <=   lut_pipe_dout_out        [(ii+1)*32-1 -: 32]       ;
//     end  


// end


// parameter CLK_PERIOD    =     6.4 ; // 156.25Mhz
// parameter CLK_1_PERIOD  =     CLK_PERIOD/64 ;

// reg clk_1 = 1'b0 ;
//  always # (CLK_1_PERIOD/2)  clk_1 = ~clk_1 ; // 64*100Mhz

// reg [7:0] seg_cnt = SEG_NUM-1 ; //  在这里8字节为一段，一拍（beat）传输64段(模拟总线位宽4096bits)



// always @( posedge clk_1 ) begin

//         if ( seg_cnt == SEG_NUM-1 )
//             seg_cnt <= 0 ;
//         else 
//             seg_cnt <=seg_cnt+1'b1 ;    

// end



// reg              seri_eop_out        ='b0   ;
// reg              seri_dval_out       ='b0   ;
// reg  [3:0]       seri_packet_num_out ='b0   ;
// reg  [31:0]      seri_dout_out       ='b0   ;


// wire [7:0] seg_cnt_process ;

// assign seg_cnt_process = ( seg_cnt>30 )?(94-seg_cnt):(30-seg_cnt) ;


// always @( posedge clk_1 ) begin
//         seri_eop_out        <= seri_lut_pipe_eop_out        [seg_cnt_process] ;
//         seri_dval_out       <= seri_lut_pipe_dval_out       [seg_cnt_process] ;
//         seri_packet_num_out <= seri_lut_pipe_packet_num_out [seg_cnt_process] ;
//         seri_dout_out       <= seri_lut_pipe_dout_out       [seg_cnt_process] ;
// end

// reg seri_eop_out_ff ;

// always @( posedge clk_1 ) begin
//     seri_eop_out_ff <= seri_eop_out ;
// end

// reg [31:0]  pkt_1_resault = 'b0  ;
// reg [31:0]  pkt_2_resault = 'b0  ;
// reg [31:0]  pkt_3_resault = 'b0  ;
// reg [31:0]  pkt_4_resault = 'b0  ;
// reg [31:0]  pkt_5_resault = 'b0  ;
// reg [31:0]  pkt_6_resault = 'b0  ;
// reg [31:0]  pkt_7_resault = 'b0  ;
// reg [31:0]  pkt_8_resault = 'b0  ;

// always @( posedge clk_1 ) begin
//     if ( seri_eop_out_ff ) begin
//         pkt_1_resault <= 'b0 ;
//     end
//     else if ( seri_dval_out == 1'b1 && seri_packet_num_out == 'd1 ) begin
//         pkt_1_resault <= pkt_1_resault ^ seri_dout_out ;
//     end
//     else begin
//         pkt_1_resault <= pkt_1_resault ;
//     end
// end

// always @( posedge clk_1 ) begin
//     if ( seri_eop_out_ff ) begin
//         pkt_2_resault <= 'b0 ;
//     end
//     else if ( seri_dval_out == 1'b1 && seri_packet_num_out == 'd2 ) begin
//         pkt_2_resault <= pkt_2_resault ^ seri_dout_out ;
//     end
//     else begin
//         pkt_2_resault <= pkt_2_resault ;
//     end
// end

// always @( posedge clk_1 ) begin
//     if ( seri_eop_out_ff ) begin
//         pkt_3_resault <= 'b0 ;
//     end
//     else if ( seri_dval_out == 1'b1 && seri_packet_num_out == 'd3 ) begin
//         pkt_3_resault <= pkt_3_resault ^ seri_dout_out ;
//     end
//     else begin
//         pkt_3_resault <= pkt_3_resault ;
//     end
// end

// always @( posedge clk_1 ) begin
//     if ( seri_eop_out_ff ) begin
//         pkt_4_resault <= 'b0 ;
//     end
//     else if ( seri_dval_out == 1'b1 && seri_packet_num_out == 'd4 ) begin
//         pkt_4_resault <= pkt_4_resault ^ seri_dout_out ;
//     end
//     else begin
//         pkt_4_resault <= pkt_4_resault ;
//     end
// end

// always @( posedge clk_1) begin
//     if ( seri_eop_out_ff ) begin
//         pkt_5_resault <= 'b0 ;
//     end
//     else if ( seri_dval_out == 1'b1 && seri_packet_num_out == 'd5 ) begin
//         pkt_5_resault <= pkt_5_resault ^ seri_dout_out ;
//     end
//     else begin
//         pkt_5_resault <= pkt_5_resault ;
//     end
// end

// always @( posedge clk_1 ) begin
//     if ( seri_eop_out_ff ) begin
//         pkt_6_resault <= 'b0 ;
//     end
//     else if ( seri_dval_out == 1'b1 && seri_packet_num_out == 'd6 ) begin
//         pkt_6_resault <= pkt_6_resault ^ seri_dout_out ;
//     end
//     else begin
//         pkt_6_resault <= pkt_6_resault ;
//     end
// end

// always @( posedge clk_1 ) begin
//     if ( seri_eop_out_ff ) begin
//         pkt_7_resault <= 'b0 ;
//     end
//     else if ( seri_dval_out == 1'b1 && seri_packet_num_out == 'd7 ) begin
//         pkt_7_resault <= pkt_7_resault ^ seri_dout_out ;
//     end
//     else begin
//         pkt_7_resault <= pkt_7_resault ;
//     end
// end

// always @( posedge clk_1 ) begin
//     if ( seri_eop_out_ff ) begin
//         pkt_8_resault <= 'b0 ;
//     end
//     else if ( seri_dval_out == 1'b1 && seri_packet_num_out == 'd8 ) begin
//         pkt_8_resault <= pkt_8_resault ^ seri_dout_out ;
//     end
//     else begin
//         pkt_8_resault <= pkt_8_resault ;
//     end
// end




//*********************
endmodule   






// 

// wire                dval_c_xor  ;
// wire [MOD_WIDTH-1:0]   mod_c_xor  ;
// wire [31:0]         dout_c_xor  ;


//  c_xor_lut_top 

// # (    .MOD_WIDTH ( MOD_WIDTH )
  
   

//   ) u_c_xor_lut_top
// ( 
//             .clk     ( clk )  ,
//             .rst     ( rst )  ,
//             .eop_in  (   )  ,
//             .dval_in (  )  ,
//             .mod_in  (   )  ,
//             .din     (  )  ,
//             .mod_out ( mod_c_xor )  ,
//             .cout_en ( dval_c_xor )  ,
//             .cout    ( dout_c_xor )  


//  ) ;






//   go_back_pipe 

// # (     
//                 .GO_BACK_STAGE( GO_BACK_STAGE    ) ,
//                 .BUS_WIDTH    ( BUS_WIDTH  ) ,
//                 .MOD_WIDTH    ( MOD_WIDTH  ) 

// ) u_go_back_pipe

//   (     
//             .clk         ( clk        )  ,
//             .rst         ( rst        )  ,
//             .crc_in      ( dout_c_xor )  ,
//             .crc_en_in   ( dval_c_xor )  ,
//             .mod_in      ( mod_c_xor  )  ,
//             .crc_out     ( crc_pre    )  ,
//             .crc_out_en  ( crc_en_pre )      
//                ) ;