
// **************************************************************
// COPYRIGHT(c)2015, Xidian University
// All rights reserved.
//
// IP LIB INDEX :  
// IP Name      :      
// File name    : 
// Module name  : 
// Full name    :  
//
// Author       : Liu-Huan 
// Email        : assasin9997@163.com 
// Data         : 
// Version      : V 1.0 
// 
// Abstract     : 
// Called by    :  
// 
// Modification history
// -----------------------------------------------------------------
// 
// 
//
// *****************************************************************

// *******************
// TIMESCALE
// ******************* 
`timescale 1ns/1ps 

// *******************
// INFORMATION
// *******************


//*******************
//DEFINE(s)
//*******************
//`define UDLY 1    //Unit delay, for non-blocking assignments in sequential logic


//*******************
//DEFINE MODULE PORT
//*******************
module  data_source_64   (     
            input 				clk     ,
            output  			sop     ,
            output  			eop     ,
            output  			dval    ,
            output  [2:0] 		mod     ,
            output  [63:0] 		dout         
              ) ;

//*******************
//DEFINE LOCAL PARAMETER
//*******************
//parameter(s)
                                    
 

//*********************
//INNER SIGNAL DECLARATION
//*********************
//REGS
  reg [79:0] mem [0:8191] ;
  reg [79:0] dout_ff = 80'b0 ;

//WIRES
 

//*********************
//INSTANTCE MODULE
//*********************

initial begin
mem[0]    = 80'h00000000000000000000;
mem[1]    = 80'h00000000000000000000;
mem[2]    = 80'h10100000010000010010;
mem[3]    = 80'h00109400000208004500;
mem[4]    = 80'h0010002e28e30000fffd;
mem[5]    = 80'h00101097c0550102c000;
mem[6]    = 80'h00100001ffabffabffab;
mem[7]    = 80'h00101c9312ab44b71a18;
mem[8]    = 80'h00103894babc2edacd5b;
mem[9]    = 80'h011026ab5bc0c1b9d9ab;
mem[10]   = 80'h00000000000000000000;
mem[11]   = 80'h10100000010000010010;
mem[12]   = 80'h00109400000208004500;
mem[13]   = 80'h0010002e28e40000fffd;
mem[14]   = 80'h00101096c0550102c000;
mem[15]   = 80'h00100001ffabffabffab;
mem[16]   = 80'h00101bb7d64195a39598;
mem[17]   = 80'h0010807babd0123becbe;
mem[18]   = 80'h011056236161ad8a4a35;
mem[19]   = 80'h00000000000000000000;
mem[20]   = 80'h00000000000000000000;
mem[21]   = 80'h00000000000000000000;
mem[22]   = 80'h10100000010000010010;
mem[23]   = 80'h00109400000208004500;
mem[24]   = 80'h0010002e28e50000fffd;
mem[25]   = 80'h00101095c0550102c000;
mem[26]   = 80'h00100001ffabffabffab;
mem[27]   = 80'h00101ac6086d4dda5727;
mem[28]   = 80'h00104ba92c3de7ebadef;
mem[29]   = 80'h0110191410f5a4d1c777;
mem[30]   = 80'h00000000000000000000;
mem[31]   = 80'h10100000010000010010;
mem[32]   = 80'h00109400000208004500;
mem[33]   = 80'h0010002e28e60000fffd;
mem[34]   = 80'h00101094c0550102c000;
mem[35]   = 80'h00100001ffabffabffab;
mem[36]   = 80'h001019546a18255010e7;
mem[37]   = 80'h001017dea40bf9a4e81d;
mem[38]   = 80'h011080c627e95b83d31b;
mem[39]   = 80'h00000000000000000000;
mem[40]   = 80'h00000000000000000000;
mem[41]   = 80'h00000000000000000000;
mem[42]   = 80'h10100000010000010010;
mem[43]   = 80'h00109400000208004500;
mem[44]   = 80'h0010002e28e70000fffd;
mem[45]   = 80'h00101093c0550102c000;
mem[46]   = 80'h00100001ffabffabffab;
mem[47]   = 80'h00101825b434fd29d258;
mem[48]   = 80'h0010dc0c23e60c74914c;
mem[49]   = 80'h011043cd82a219d42b40;
mem[50]   = 80'h00000000000000000000;
mem[51]   = 80'h10100000010000010010;
mem[52]   = 80'h00109400000208004500;
mem[53]   = 80'h0010002e28e80000fffd;
mem[54]   = 80'h00101092c0550102c000;
mem[55]   = 80'h00100001ffabffabffab;
mem[56]   = 80'h0010171de3cd87790fe6;
mem[57]   = 80'h0010660086d380666dd6;
mem[58]   = 80'h0110cd05c59e6c633f86;
mem[59]   = 80'h00000000000000000000;
mem[60]   = 80'h00000000000000000000;
mem[61]   = 80'h00000000000000000000;
mem[62]   = 80'h10100000010000010010;
mem[63]   = 80'h00109400000208004500;
mem[64]   = 80'h0010002e28e90000fffd;
mem[65]   = 80'h00101091c0550102c000;
mem[66]   = 80'h00100001ffabffabffab;
mem[67]   = 80'h0010166c3de15f00cd59;
mem[68]   = 80'h0010add2013e75b66487;
mem[69]   = 80'h01100657efb2e2276b97;
mem[70]   = 80'h00000000000000000000;
mem[71]   = 80'h00000000000000000000;
mem[72]   = 80'h00000000000000000000;
mem[73]   = 80'h10100000010000010010;
mem[74]   = 80'h00109400000208004500;
mem[75]   = 80'h0010002e28ea0000fffd;
mem[76]   = 80'h00101090c0550102c000;
mem[77]   = 80'h00100001ffabffabffab;
mem[78]   = 80'h001015fe5f94378a8a99;
mem[79]   = 80'h0010f1a589086bc6f175;
mem[80]   = 80'h011063368d28dbdad57f;
mem[81]   = 80'h00000000000000000000;
mem[82]   = 80'h00000000000000000000;
mem[83]   = 80'h00000000000000000000;
mem[84]   = 80'h10100000010000010010;
mem[85]   = 80'h00109400000208004500;
mem[86]   = 80'h0010002e28eb0000fffd;
mem[87]   = 80'h0010108fc0550102c000;
mem[88]   = 80'h00100001ffabffabffab;
mem[89]   = 80'h0010148f81b8eff34826;
mem[90]   = 80'h00103a770ee59e167324;
mem[91]   = 80'h01106f066800cb0a15fc;
mem[92]   = 80'h00000000000000000000;
mem[93]   = 80'h10100000010000010010;
mem[94]   = 80'h00109400000208004500;
mem[95]   = 80'h0010002e28ec0000fffd;
mem[96]   = 80'h0010108ec0550102c000;
mem[97]   = 80'h00100001ffabffabffab;
mem[98]   = 80'h001013ab45523ee7c7a6;
mem[99]   = 80'h001082981f89a2f701c1;
mem[100]  = 80'h011044621538bb108362;
mem[101]  = 80'h00000000000000000000;
mem[102]  = 80'h00000000000000000000;
mem[103]  = 80'h00000000000000000000;
mem[104]  = 80'h00000000000000000000;
mem[105]  = 80'h10100000010000010010;
mem[106]  = 80'h00109400000208004500;
mem[107]  = 80'h0010002e28ed0000fffd;
mem[108]  = 80'h0010108dc0550102c000;
mem[109]  = 80'h00100001ffabffabffab;
mem[110]  = 80'h001012da9b7ee69e0519;
mem[111]  = 80'h0010494a986457277f90;
mem[112]  = 80'h01101efe8e8a7d755411;
mem[113]  = 80'h00000000000000000000;
mem[114]  = 80'h00000000000000000000;
mem[115]  = 80'h00000000000000000000;
mem[116]  = 80'h10100000010000010010;
mem[117]  = 80'h00109400000208004500;
mem[118]  = 80'h0010002e28ee0000fffd;
mem[119]  = 80'h0010108cc0550102c000;
mem[120]  = 80'h00100001ffabffabffab;
mem[121]  = 80'h00101148f90b8e1442d9;
mem[122]  = 80'h0010153d10524957b662;
mem[123]  = 80'h0110304dcf27c4acaa46;
mem[124]  = 80'h00000000000000000000;
mem[125]  = 80'h10100000010000010010;
mem[126]  = 80'h00109400000208004500;
mem[127]  = 80'h0010002e28ef0000fffd;
mem[128]  = 80'h0010108bc0550102c000;
mem[129]  = 80'h00100001ffabffabffab;
mem[130]  = 80'h001010392727566d8066;
mem[131]  = 80'h0010deef97bfbc87ff33;
mem[132]  = 80'h0110f6d3c88c114a15e9;
mem[133]  = 80'h00000000000000000000;
mem[134]  = 80'h00000000000000000000;
mem[135]  = 80'h00000000000000000000;
mem[136]  = 80'h00000000000000000000;
mem[137]  = 80'h10100000010000010010;
mem[138]  = 80'h00109400000208004500;
mem[139]  = 80'h0010002e28f00000fffd;
mem[140]  = 80'h0010108ac0550102c000;
mem[141]  = 80'h00100001ffabffabffab;
mem[142]  = 80'h00100f3856f97ab5f9a4;
mem[143]  = 80'h001061245a395173cb56;
mem[144]  = 80'h0110dd906fbb2c1df4f8;
mem[145]  = 80'h00000000000000000000;
mem[146]  = 80'h00000000000000000000;
mem[147]  = 80'h00000000000000000000;
mem[148]  = 80'h10100000010000010010;
mem[149]  = 80'h00109400000208004500;
mem[150]  = 80'h0010002e28f10000fffd;
mem[151]  = 80'h00101089c0550102c000;
mem[152]  = 80'h00100001ffabffabffab;
mem[153]  = 80'h00100e4988d5a2cc3b1b;
mem[154]  = 80'h0010aaf6ddd4a4a39407;
mem[155]  = 80'h0110b2db16a7de9ac655;
mem[156]  = 80'h00000000000000000000;
mem[157]  = 80'h10100000010000010010;
mem[158]  = 80'h00109400000208004500;
mem[159]  = 80'h0010002e28f20000fffd;
mem[160]  = 80'h00101088c0550102c000;
mem[161]  = 80'h00100001ffabffabffab;
mem[162]  = 80'h00100ddbeaa0ca467cdb;
mem[163]  = 80'h0010f68155e2bad357f5;
mem[164]  = 80'h011073a3ed90a674b5be;
mem[165]  = 80'h00000000000000000000;
mem[166]  = 80'h00000000000000000000;
mem[167]  = 80'h00000000000000000000;
mem[168]  = 80'h10100000010000010010;
mem[169]  = 80'h00109400000208004500;
mem[170]  = 80'h0010002e28f30000fffd;
mem[171]  = 80'h00101087c0550102c000;
mem[172]  = 80'h00100001ffabffabffab;
mem[173]  = 80'h00100caa348c123fbe64;
mem[174]  = 80'h00103d53d20f4f0314a4;
mem[175]  = 80'h01105af62025783a28a2;
mem[176]  = 80'h00000000000000000000;
mem[177]  = 80'h00000000000000000000;
mem[178]  = 80'h00000000000000000000;
mem[179]  = 80'h10100000010000010010;
mem[180]  = 80'h00109400000208004500;
mem[181]  = 80'h0010002e28f40000fffd;
mem[182]  = 80'h00101086c0550102c000;
mem[183]  = 80'h00100001ffabffabffab;
mem[184]  = 80'h00100b8ef066c32b31e4;
mem[185]  = 80'h001085bcc36373e25641;
mem[186]  = 80'h0110740787afb9527aaa;
mem[187]  = 80'h00000000000000000000;
mem[188]  = 80'h00000000000000000000;
mem[189]  = 80'h00000000000000000000;
mem[190]  = 80'h10100000010000010010;
mem[191]  = 80'h00109400000208004500;
mem[192]  = 80'h0010002e28f50000fffd;
mem[193]  = 80'h00101085c0550102c000;
mem[194]  = 80'h00100001ffabffabffab;
mem[195]  = 80'h00100aff2e4a1b52f35b;
mem[196]  = 80'h00104e6e448e8632d810;
mem[197]  = 80'h01103d5a896eb974c4db;
mem[198]  = 80'h00000000000000000000;
mem[199]  = 80'h10100000010000010010;
mem[200]  = 80'h00109400000208004500;
mem[201]  = 80'h0010002e28f60000fffd;
mem[202]  = 80'h00101084c0550102c000;
mem[203]  = 80'h00100001ffabffabffab;
mem[204]  = 80'h0010096d4c3f73d8b49b;
mem[205]  = 80'h00101219ccb8984252e2;
mem[206]  = 80'h01104b766c72b5f70d8b;
mem[207]  = 80'h00000000000000000000;
mem[208]  = 80'h00000000000000000000;
mem[209]  = 80'h00000000000000000000;
mem[210]  = 80'h10100000010000010010;
mem[211]  = 80'h00109400000208004500;
mem[212]  = 80'h0010002e28f70000fffd;
mem[213]  = 80'h00101083c0550102c000;
mem[214]  = 80'h00100001ffabffabffab;
mem[215]  = 80'h0010081c9213aba17624;
mem[216]  = 80'h0010d9cb4b556d9249b3;
mem[217]  = 80'h0110e535826d23fe875d;
mem[218]  = 80'h00000000000000000000;
mem[219]  = 80'h00000000000000000000;
mem[220]  = 80'h00000000000000000000;
mem[221]  = 80'h10100000010000010010;
mem[222]  = 80'h00109400000208004500;
mem[223]  = 80'h0010002e28f80000fffd;
mem[224]  = 80'h00101082c0550102c000;
mem[225]  = 80'h00100001ffabffabffab;
mem[226]  = 80'h00100724c5ead1f1ab9a;
mem[227]  = 80'h001063c7ee60e180b729;
mem[228]  = 80'h01100d9fbcf2216f6732;
mem[229]  = 80'h00000000000000000000;
mem[230]  = 80'h00000000000000000000;
mem[231]  = 80'h00000000000000000000;
mem[232]  = 80'h10100000010000010010;
mem[233]  = 80'h00109400000208004500;
mem[234]  = 80'h0010002e28f90000fffd;
mem[235]  = 80'h00101081c0550102c000;
mem[236]  = 80'h00100001ffabffabffab;
mem[237]  = 80'h001006551bc609886925;
mem[238]  = 80'h0010a815698d14533878;
mem[239]  = 80'h01102ea3de2593a77f99;
mem[240]  = 80'h00000000000000000000;
mem[241]  = 80'h10100000010000010010;
mem[242]  = 80'h00109400000208004500;
mem[243]  = 80'h0010002e28fa0000fffd;
mem[244]  = 80'h00101080c0550102c000;
mem[245]  = 80'h00100001ffabffabffab;
mem[246]  = 80'h001005c779b361022ee5;
mem[247]  = 80'h0010f462e1bb0a238b8a;
mem[248]  = 80'h0110e7829d4e95403691;
mem[249]  = 80'h00000000000000000000;
mem[250]  = 80'h00000000000000000000;
mem[251]  = 80'h00000000000000000000;
mem[252]  = 80'h00000000000000000000;
mem[253]  = 80'h10100000010000010010;
mem[254]  = 80'h00109400000208004500;
mem[255]  = 80'h0010002e28fb0000fffd;
mem[256]  = 80'h0010107fc0550102c000;
mem[257]  = 80'h00100001ffabffabffab;
mem[258]  = 80'h001004b6a79fb97bec5a;
mem[259]  = 80'h00103fb06656fff3cadb;
mem[260]  = 80'h0110a8b594471706ebde;
mem[261]  = 80'h00000000000000000000;
mem[262]  = 80'h00000000000000000000;
mem[263]  = 80'h00000000000000000000;
mem[264]  = 80'h10100000010000010010;
mem[265]  = 80'h00109400000208004500;
mem[266]  = 80'h0010002e28fc0000fffd;
mem[267]  = 80'h0010107ec0550102c000;
mem[268]  = 80'h00100001ffabffabffab;
mem[269]  = 80'h001003926375686f63da;
mem[270]  = 80'h0010875f773ac312fb3e;
mem[271]  = 80'h0110db4e3474ffde0392;
mem[272]  = 80'h00000000000000000000;
mem[273]  = 80'h10100000010000010010;
mem[274]  = 80'h00109400000208004500;
mem[275]  = 80'h0010002e28fd0000fffd;
mem[276]  = 80'h0010107dc0550102c000;
mem[277]  = 80'h00100001ffabffabffab;
mem[278]  = 80'h001002e3bd59b016a165;
mem[279]  = 80'h00104c8df0d736c2ba6f;
mem[280]  = 80'h011094792b363eb44044;
mem[281]  = 80'h00000000000000000000;
mem[282]  = 80'h00000000000000000000;
mem[283]  = 80'h00000000000000000000;
mem[284]  = 80'h10100000010000010010;
mem[285]  = 80'h00109400000208004500;
mem[286]  = 80'h0010002e28fe0000fffd;
mem[287]  = 80'h0010107cc0550102c000;
mem[288]  = 80'h00100001ffabffabffab;
mem[289]  = 80'h00100171df2cd89ce6a5;
mem[290]  = 80'h001010fa78e128b2ef9d;
mem[291]  = 80'h0110e74cd6a657a6ddb5;
mem[292]  = 80'h00000000000000000000;
mem[293]  = 80'h10100000010000010010;
mem[294]  = 80'h00109400000208004500;
mem[295]  = 80'h0010002e28ff0000fffd;
mem[296]  = 80'h0010107bc0550102c000;
mem[297]  = 80'h00100001ffabffabffab;
mem[298]  = 80'h00100000010000e5241a;
mem[299]  = 80'h0010db28ff0cdd62a5cc;
mem[300]  = 80'h01107481081ac4a6f6dd;
mem[301]  = 80'h00000000000000000000;
mem[302]  = 80'h00000000000000000000;
mem[303]  = 80'h00000000000000000000;
mem[304]  = 80'h00000000000000000000;
mem[305]  = 80'h10100000010000010010;
mem[306]  = 80'h00109400000208004500;
mem[307]  = 80'h0010002e29000000fffd;
mem[308]  = 80'h0010107ac0550102c000;
mem[309]  = 80'h00100001ffabffabffab;
mem[310]  = 80'h0010ff2f4b1bb732658f;
mem[311]  = 80'h00109d9882578e2d1c03;
mem[312]  = 80'h0110234dab84cb920ef7;
mem[313]  = 80'h00000000000000000000;
mem[314]  = 80'h00000000000000000000;
mem[315]  = 80'h00000000000000000000;
mem[316]  = 80'h10100000010000010010;
mem[317]  = 80'h00109400000208004500;
mem[318]  = 80'h0010002e29010000fffd;
mem[319]  = 80'h00101079c0550102c000;
mem[320]  = 80'h00100001ffabffabffab;
mem[321]  = 80'h0010fe5e95376f4ba730;
mem[322]  = 80'h0010564a05ba7bfd6252;
mem[323]  = 80'h011079d1a1c7dc8e3926;
mem[324]  = 80'h00000000000000000000;
mem[325]  = 80'h00000000000000000000;
mem[326]  = 80'h00000000000000000000;
mem[327]  = 80'h10100000010000010010;
mem[328]  = 80'h00109400000208004500;
mem[329]  = 80'h0010002e29020000fffd;
mem[330]  = 80'h00101078c0550102c000;
mem[331]  = 80'h00100001ffabffabffab;
mem[332]  = 80'h0010fdccf74207c1e0f0;
mem[333]  = 80'h00100a3d8d8c658de3a0;
mem[334]  = 80'h0110d3076e3eebd7ed77;
mem[335]  = 80'h00000000000000000000;
mem[336]  = 80'h10100000010000010010;
mem[337]  = 80'h00109400000208004500;
mem[338]  = 80'h0010002e29030000fffd;
mem[339]  = 80'h00101077c0550102c000;
mem[340]  = 80'h00100001ffabffabffab;
mem[341]  = 80'h0010fcbd296edfb8224f;
mem[342]  = 80'h0010c1ef0a61905c62f1;
mem[343]  = 80'h0110bd545ad8b26b75a4;
mem[344]  = 80'h00000000000000000000;
mem[345]  = 80'h00000000000000000000;
mem[346]  = 80'h00000000000000000000;
mem[347]  = 80'h10100000010000010010;
mem[348]  = 80'h00109400000208004500;
mem[349]  = 80'h0010002e29040000fffd;
mem[350]  = 80'h00101076c0550102c000;
mem[351]  = 80'h00100001ffabffabffab;
mem[352]  = 80'h0010fb99ed840eacadcf;
mem[353]  = 80'h001079001b0dacbd0714;
mem[354]  = 80'h01100cd405b2a54cf17a;
mem[355]  = 80'h00000000000000000000;
mem[356]  = 80'h10100000010000010010;
mem[357]  = 80'h00109400000208004500;
mem[358]  = 80'h0010002e29050000fffd;
mem[359]  = 80'h00101075c0550102c000;
mem[360]  = 80'h00100001ffabffabffab;
mem[361]  = 80'h0010fae833a8d6d56f70;
mem[362]  = 80'h0010b2d29ce0596d0e45;
mem[363]  = 80'h0110c7860c3c8ebdd4ed;
mem[364]  = 80'h00000000000000000000;
mem[365]  = 80'h00000000000000000000;
mem[366]  = 80'h00000000000000000000;
mem[367]  = 80'h00000000000000000000;
mem[368]  = 80'h10100000010000010010;
mem[369]  = 80'h00109400000208004500;
mem[370]  = 80'h0010002e29060000fffd;
mem[371]  = 80'h00101074c0550102c000;
mem[372]  = 80'h00100001ffabffabffab;
mem[373]  = 80'h0010f97a51ddbe5f28b0;
mem[374]  = 80'h0010eea514d6471d87b7;
mem[375]  = 80'h0110e4f9164dc2c38709;
mem[376]  = 80'h00000000000000000000;
mem[377]  = 80'h00000000000000000000;
mem[378]  = 80'h00000000000000000000;
mem[379]  = 80'h10100000010000010010;
mem[380]  = 80'h00109400000208004500;
mem[381]  = 80'h0010002e29070000fffd;
mem[382]  = 80'h00101073c0550102c000;
mem[383]  = 80'h00100001ffabffabffab;
mem[384]  = 80'h0010f80b8ff16626ea0f;
mem[385]  = 80'h00102577933bb2cdfee6;
mem[386]  = 80'h011027f2957281a2c9c6;
mem[387]  = 80'h00000000000000000000;
mem[388]  = 80'h00000000000000000000;
mem[389]  = 80'h00000000000000000000;
mem[390]  = 80'h10100000010000010010;
mem[391]  = 80'h00109400000208004500;
mem[392]  = 80'h0010002e29080000fffd;
mem[393]  = 80'h00101072c0550102c000;
mem[394]  = 80'h00100001ffabffabffab;
mem[395]  = 80'h0010f733d8081c7637b1;
mem[396]  = 80'h00109f7b360e3edfc07c;
mem[397]  = 80'h0110d90c2ea99f4a4391;
mem[398]  = 80'h00000000000000000000;
mem[399]  = 80'h10100000010000010010;
mem[400]  = 80'h00109400000208004500;
mem[401]  = 80'h0010002e29090000fffd;
mem[402]  = 80'h00101071c0550102c000;
mem[403]  = 80'h00100001ffabffabffab;
mem[404]  = 80'h0010f6420624c40ff50e;
mem[405]  = 80'h001054a9b1e3cb0f8f2d;
mem[406]  = 80'h0110b534347bc261a949;
mem[407]  = 80'h00000000000000000000;
mem[408]  = 80'h00000000000000000000;
mem[409]  = 80'h00000000000000000000;
mem[410]  = 80'h00000000000000000000;
mem[411]  = 80'h10100000010000010010;
mem[412]  = 80'h00109400000208004500;
mem[413]  = 80'h0010002e290a0000fffd;
mem[414]  = 80'h00101070c0550102c000;
mem[415]  = 80'h00100001ffabffabffab;
mem[416]  = 80'h0010f5d06451ac85b2ce;
mem[417]  = 80'h001008de39d5d57f5ddf;
mem[418]  = 80'h0110440e8c689c07320e;
mem[419]  = 80'h00000000000000000000;
mem[420]  = 80'h00000000000000000000;
mem[421]  = 80'h00000000000000000000;
mem[422]  = 80'h10100000010000010010;
mem[423]  = 80'h00109400000208004500;
mem[424]  = 80'h0010002e290b0000fffd;
mem[425]  = 80'h0010106fc0550102c000;
mem[426]  = 80'h00100001ffabffabffab;
mem[427]  = 80'h0010f4a1ba7d74fc7071;
mem[428]  = 80'h0010c30cbe3820af1f8e;
mem[429]  = 80'h01105e6a4b85083761ce;
mem[430]  = 80'h00000000000000000000;
mem[431]  = 80'h10100000010000010010;
mem[432]  = 80'h00109400000208004500;
mem[433]  = 80'h0010002e290c0000fffd;
mem[434]  = 80'h0010106ec0550102c000;
mem[435]  = 80'h00100001ffabffabffab;
mem[436]  = 80'h0010f3857e97a5e8fff1;
mem[437]  = 80'h00107be3af541c49ad6b;
mem[438]  = 80'h0110e6ca0c50283df946;
mem[439]  = 80'h00000000000000000000;
mem[440]  = 80'h00000000000000000000;
mem[441]  = 80'h00000000000000000000;
mem[442]  = 80'h10100000010000010010;
mem[443]  = 80'h00109400000208004500;
mem[444]  = 80'h0010002e290d0000fffd;
mem[445]  = 80'h0010106dc0550102c000;
mem[446]  = 80'h00100001ffabffabffab;
mem[447]  = 80'h0010f2f4a0bb7d913d4e;
mem[448]  = 80'h0010b03128b9e999d23a;
mem[449]  = 80'h01108f678d488ee36bbf;
mem[450]  = 80'h00000000000000000000;
mem[451]  = 80'h00000000000000000000;
mem[452]  = 80'h00000000000000000000;
mem[453]  = 80'h10100000010000010010;
mem[454]  = 80'h00109400000208004500;
mem[455]  = 80'h0010002e290e0000fffd;
mem[456]  = 80'h0010106cc0550102c000;
mem[457]  = 80'h00100001ffabffabffab;
mem[458]  = 80'h0010f166c2ce151b7a8e;
mem[459]  = 80'h0010ec46a08ff7e959c8;
mem[460]  = 80'h0110ca7a131dc6320220;
mem[461]  = 80'h00000000000000000000;
mem[462]  = 80'h00000000000000000000;
mem[463]  = 80'h00000000000000000000;
mem[464]  = 80'h10100000010000010010;
mem[465]  = 80'h00109400000208004500;
mem[466]  = 80'h0010002e290f0000fffd;
mem[467]  = 80'h0010106bc0550102c000;
mem[468]  = 80'h00100001ffabffabffab;
mem[469]  = 80'h0010f0171ce2cd62b831;
mem[470]  = 80'h00102794276202395299;
mem[471]  = 80'h0110674a625e26cb5825;
mem[472]  = 80'h00000000000000000000;
mem[473]  = 80'h10100000010000010010;
mem[474]  = 80'h00109400000208004500;
mem[475]  = 80'h0010002e29100000fffd;
mem[476]  = 80'h0010106ac0550102c000;
mem[477]  = 80'h00100001ffabffabffab;
mem[478]  = 80'h0010ef166d3ce1bac1f3;
mem[479]  = 80'h0010985feae4efcca6fc;
mem[480]  = 80'h01106d6d7882b9c9c5b2;
mem[481]  = 80'h00000000000000000000;
mem[482]  = 80'h00000000000000000000;
mem[483]  = 80'h00000000000000000000;
mem[484]  = 80'h10100000010000010010;
mem[485]  = 80'h00109400000208004500;
mem[486]  = 80'h0010002e29110000fffd;
mem[487]  = 80'h00101069c0550102c000;
mem[488]  = 80'h00100001ffabffabffab;
mem[489]  = 80'h0010ee67b31039c3034c;
mem[490]  = 80'h0010538d6d091a1c39ad;
mem[491]  = 80'h01101472f8a5006dad64;
mem[492]  = 80'h00000000000000000000;
mem[493]  = 80'h10100000010000010010;
mem[494]  = 80'h00109400000208004500;
mem[495]  = 80'h0010002e29120000fffd;
mem[496]  = 80'h00101068c0550102c000;
mem[497]  = 80'h00100001ffabffabffab;
mem[498]  = 80'h0010edf5d1655149448c;
mem[499]  = 80'h00100ffae53f046cb95f;
mem[500]  = 80'h01108d956a33aa600aeb;
mem[501]  = 80'h00000000000000000000;
mem[502]  = 80'h00000000000000000000;
mem[503]  = 80'h00000000000000000000;
mem[504]  = 80'h00000000000000000000;
mem[505]  = 80'h10100000010000010010;
mem[506]  = 80'h00109400000208004500;
mem[507]  = 80'h0010002e29130000fffd;
mem[508]  = 80'h00101067c0550102c000;
mem[509]  = 80'h00100001ffabffabffab;
mem[510]  = 80'h0010ec840f4989308633;
mem[511]  = 80'h0010c42862d2f1bcbb0e;
mem[512]  = 80'h01109a3d86c94ed187f4;
mem[513]  = 80'h00000000000000000000;
mem[514]  = 80'h00000000000000000000;
mem[515]  = 80'h00000000000000000000;
mem[516]  = 80'h10100000010000010010;
mem[517]  = 80'h00109400000208004500;
mem[518]  = 80'h0010002e29140000fffd;
mem[519]  = 80'h00101066c0550102c000;
mem[520]  = 80'h00100001ffabffabffab;
mem[521]  = 80'h0010eba0cba3582409b3;
mem[522]  = 80'h00107cc773becd5dfaeb;
mem[523]  = 80'h0110e19f4c74bd148680;
mem[524]  = 80'h00000000000000000000;
mem[525]  = 80'h00000000000000000000;
mem[526]  = 80'h00000000000000000000;
mem[527]  = 80'h10100000010000010010;
mem[528]  = 80'h00109400000208004500;
mem[529]  = 80'h0010002e29150000fffd;
mem[530]  = 80'h00101065c0550102c000;
mem[531]  = 80'h00100001ffabffabffab;
mem[532]  = 80'h0010ead1158f805dcb0c;
mem[533]  = 80'h0010b715f453388db4ba;
mem[534]  = 80'h0110be965ceca974e138;
mem[535]  = 80'h00000000000000000000;
mem[536]  = 80'h00000000000000000000;
mem[537]  = 80'h00000000000000000000;
mem[538]  = 80'h10100000010000010010;
mem[539]  = 80'h00109400000208004500;
mem[540]  = 80'h0010002e29160000fffd;
mem[541]  = 80'h00101064c0550102c000;
mem[542]  = 80'h00100001ffabffabffab;
mem[543]  = 80'h0010e94377fae8d78ccc;
mem[544]  = 80'h0010eb627c6526fcfe48;
mem[545]  = 80'h0110e9deb230795277f0;
mem[546]  = 80'h00000000000000000000;
mem[547]  = 80'h10100000010000010010;
mem[548]  = 80'h00109400000208004500;
mem[549]  = 80'h0010002e29170000fffd;
mem[550]  = 80'h00101063c0550102c000;
mem[551]  = 80'h00100001ffabffabffab;
mem[552]  = 80'h0010e832a9d630ae4e73;
mem[553]  = 80'h001020b0fb88d32ca419;
mem[554]  = 80'h01107960e1f49e367b0f;
mem[555]  = 80'h00000000000000000000;
mem[556]  = 80'h00000000000000000000;
mem[557]  = 80'h00000000000000000000;
mem[558]  = 80'h10100000010000010010;
mem[559]  = 80'h00109400000208004500;
mem[560]  = 80'h0010002e29180000fffd;
mem[561]  = 80'h00101062c0550102c000;
mem[562]  = 80'h00100001ffabffabffab;
mem[563]  = 80'h0010e70afe2f4afe93cd;
mem[564]  = 80'h00109abc5ebd5f3e1483;
mem[565]  = 80'h0110bf090fb4ce369911;
mem[566]  = 80'h00000000000000000000;
mem[567]  = 80'h00000000000000000000;
mem[568]  = 80'h00000000000000000000;
mem[569]  = 80'h10100000010000010010;
mem[570]  = 80'h00109400000208004500;
mem[571]  = 80'h0010002e29190000fffd;
mem[572]  = 80'h00101061c0550102c000;
mem[573]  = 80'h00100001ffabffabffab;
mem[574]  = 80'h0010e67b200392875172;
mem[575]  = 80'h0010516ed950aaee55d2;
mem[576]  = 80'h0110f03ef9c79014b819;
mem[577]  = 80'h00000000000000000000;
mem[578]  = 80'h10100000010000010010;
mem[579]  = 80'h00109400000208004500;
mem[580]  = 80'h0010002e291a0000fffd;
mem[581]  = 80'h00101060c0550102c000;
mem[582]  = 80'h00100001ffabffabffab;
mem[583]  = 80'h0010e5e94276fa0d16b2;
mem[584]  = 80'h00100d195166b49ee420;
mem[585]  = 80'h01105f7d702379443545;
mem[586]  = 80'h00000000000000000000;
mem[587]  = 80'h00000000000000000000;
mem[588]  = 80'h00000000000000000000;
mem[589]  = 80'h10100000010000010010;
mem[590]  = 80'h00109400000208004500;
mem[591]  = 80'h0010002e291b0000fffd;
mem[592]  = 80'h0010105fc0550102c000;
mem[593]  = 80'h00100001ffabffabffab;
mem[594]  = 80'h0010e4989c5a2274d40d;
mem[595]  = 80'h0010c6cbd68b414e6571;
mem[596]  = 80'h0110061e3e55f9189c8c;
mem[597]  = 80'h00000000000000000000;
mem[598]  = 80'h00000000000000000000;
mem[599]  = 80'h00000000000000000000;
mem[600]  = 80'h10100000010000010010;
mem[601]  = 80'h00109400000208004500;
mem[602]  = 80'h0010002e291c0000fffd;
mem[603]  = 80'h0010105ec0550102c000;
mem[604]  = 80'h00100001ffabffabffab;
mem[605]  = 80'h0010e3bc58b0f3605b8d;
mem[606]  = 80'h00107e24c7e77daf1094;
mem[607]  = 80'h0110b4edeb6603dd17c6;
mem[608]  = 80'h00000000000000000000;
mem[609]  = 80'h10100000010000010010;
mem[610]  = 80'h00109400000208004500;
mem[611]  = 80'h0010002e291d0000fffd;
mem[612]  = 80'h0010105dc0550102c000;
mem[613]  = 80'h00100001ffabffabffab;
mem[614]  = 80'h0010e2cd869c2b199932;
mem[615]  = 80'h0010b5f6400a887f08c5;
mem[616]  = 80'h01104ffdfb067e3a3fc6;
mem[617]  = 80'h00000000000000000000;
mem[618]  = 80'h00000000000000000000;
mem[619]  = 80'h00000000000000000000;
mem[620]  = 80'h00000000000000000000;
mem[621]  = 80'h10100000010000010010;
mem[622]  = 80'h00109400000208004500;
mem[623]  = 80'h0010002e291e0000fffd;
mem[624]  = 80'h0010105cc0550102c000;
mem[625]  = 80'h00100001ffabffabffab;
mem[626]  = 80'h0010e15fe4e94393def2;
mem[627]  = 80'h0010e981c83c960f8037;
mem[628]  = 80'h01105fb3ef76675283c7;
mem[629]  = 80'h00000000000000000000;
mem[630]  = 80'h00000000000000000000;
mem[631]  = 80'h00000000000000000000;
mem[632]  = 80'h10100000010000010010;
mem[633]  = 80'h00109400000208004500;
mem[634]  = 80'h0010002e291f0000fffd;
mem[635]  = 80'h0010105bc0550102c000;
mem[636]  = 80'h00100001ffabffabffab;
mem[637]  = 80'h0010e02e3ac59bea1c4d;
mem[638]  = 80'h001022534fd163dc0966;
mem[639]  = 80'h0110d6297743ba782c6d;
mem[640]  = 80'h00000000000000000000;
mem[641]  = 80'h10100000010000010010;
mem[642]  = 80'h00109400000208004500;
mem[643]  = 80'h0010002e29200000fffd;
mem[644]  = 80'h0010105ac0550102c000;
mem[645]  = 80'h00100001ffabffabffab;
mem[646]  = 80'h0010df5d07551a232d77;
mem[647]  = 80'h0010961653314de7e9fd;
mem[648]  = 80'h01103a047681295bf20f;
mem[649]  = 80'h00000000000000000000;
mem[650]  = 80'h00000000000000000000;
mem[651]  = 80'h00000000000000000000;
mem[652]  = 80'h00000000000000000000;
mem[653]  = 80'h10100000010000010010;
mem[654]  = 80'h00109400000208004500;
mem[655]  = 80'h0010002e29210000fffd;
mem[656]  = 80'h00101059c0550102c000;
mem[657]  = 80'h00100001ffabffabffab;
mem[658]  = 80'h0010de2cd979c25aefc8;
mem[659]  = 80'h00105dc4d4dcb83797ac;
mem[660]  = 80'h01106098b317e4aa1e64;
mem[661]  = 80'h00000000000000000000;
mem[662]  = 80'h10100000010000010010;
mem[663]  = 80'h00109400000208004500;
mem[664]  = 80'h0010002e29220000fffd;
mem[665]  = 80'h00101058c0550102c000;
mem[666]  = 80'h00100001ffabffabffab;
mem[667]  = 80'h0010ddbebb0caad0a808;
mem[668]  = 80'h001001b35ceaa647555e;
mem[669]  = 80'h011092d12746d4fcb2c5;
mem[670]  = 80'h00000000000000000000;
mem[671]  = 80'h00000000000000000000;
mem[672]  = 80'h00000000000000000000;
mem[673]  = 80'h00000000000000000000;
mem[674]  = 80'h10100000010000010010;
mem[675]  = 80'h00109400000208004500;
mem[676]  = 80'h0010002e29230000fffd;
mem[677]  = 80'h00101057c0550102c000;
mem[678]  = 80'h00100001ffabffabffab;
mem[679]  = 80'h0010dccf652072a96ab7;
mem[680]  = 80'h0010ca61db075397160f;
mem[681]  = 80'h0110bb84161a6746f0b8;
mem[682]  = 80'h00000000000000000000;
mem[683]  = 80'h00000000000000000000;
mem[684]  = 80'h00000000000000000000;
mem[685]  = 80'h10100000010000010010;
mem[686]  = 80'h00109400000208004500;
mem[687]  = 80'h0010002e29240000fffd;
mem[688]  = 80'h00101056c0550102c000;
mem[689]  = 80'h00100001ffabffabffab;
mem[690]  = 80'h0010dbeba1caa3bde537;
mem[691]  = 80'h0010728eca6b6f76b5ea;
mem[692]  = 80'h0110b6f6e0014f8ce618;
mem[693]  = 80'h00000000000000000000;
mem[694]  = 80'h10100000010000010010;
mem[695]  = 80'h00109400000208004500;
mem[696]  = 80'h0010002e29250000fffd;
mem[697]  = 80'h00101055c0550102c000;
mem[698]  = 80'h00100001ffabffabffab;
mem[699]  = 80'h0010da9a7fe67bc42788;
mem[700]  = 80'h0010b95c4d869aa6fabb;
mem[701]  = 80'h0110dace8b1d1200f48a;
mem[702]  = 80'h00000000000000000000;
mem[703]  = 80'h00000000000000000000;
mem[704]  = 80'h00000000000000000000;
mem[705]  = 80'h00000000000000000000;
mem[706]  = 80'h10100000010000010010;
mem[707]  = 80'h00109400000208004500;
mem[708]  = 80'h0010002e29260000fffd;
mem[709]  = 80'h00101054c0550102c000;
mem[710]  = 80'h00100001ffabffabffab;
mem[711]  = 80'h0010d9081d93134e6048;
mem[712]  = 80'h0010e52bc5b084d63149;
mem[713]  = 80'h0110921fa2b1081eff1f;
mem[714]  = 80'h00000000000000000000;
mem[715]  = 80'h10100000010000010010;
mem[716]  = 80'h00109400000208004500;
mem[717]  = 80'h0010002e29270000fffd;
mem[718]  = 80'h00101053c0550102c000;
mem[719]  = 80'h00100001ffabffabffab;
mem[720]  = 80'h0010d879c3bfcb37a2f7;
mem[721]  = 80'h00102ef9425d71064a18;
mem[722]  = 80'h0110377691ab2e13a667;
mem[723]  = 80'h00000000000000000000;
mem[724]  = 80'h00000000000000000000;
mem[725]  = 80'h00000000000000000000;
mem[726]  = 80'h00000000000000000000;
mem[727]  = 80'h10100000010000010010;
mem[728]  = 80'h00109400000208004500;
mem[729]  = 80'h0010002e29280000fffd;
mem[730]  = 80'h00101052c0550102c000;
mem[731]  = 80'h00100001ffabffabffab;
mem[732]  = 80'h0010d7419446b1677f49;
mem[733]  = 80'h001094f5e768fd14bb82;
mem[734]  = 80'h0110cfe25eed70155475;
mem[735]  = 80'h00000000000000000000;
mem[736]  = 80'h10100000010000010010;
mem[737]  = 80'h00109400000208004500;
mem[738]  = 80'h0010002e29290000fffd;
mem[739]  = 80'h00101051c0550102c000;
mem[740]  = 80'h00100001ffabffabffab;
mem[741]  = 80'h0010d6304a6a691ebdf6;
mem[742]  = 80'h00105f27608508c53bd3;
mem[743]  = 80'h01109280218abb754a61;
mem[744]  = 80'h00000000000000000000;
mem[745]  = 80'h00000000000000000000;
mem[746]  = 80'h00000000000000000000;
mem[747]  = 80'h00000000000000000000;
mem[748]  = 80'h10100000010000010010;
mem[749]  = 80'h00109400000208004500;
mem[750]  = 80'h0010002e292a0000fffd;
mem[751]  = 80'h00101050c0550102c000;
mem[752]  = 80'h00100001ffabffabffab;
mem[753]  = 80'h0010d5a2281f0194fa36;
mem[754]  = 80'h00100350e8b316b5ab21;
mem[755]  = 80'h01100814508434b8be22;
mem[756]  = 80'h00000000000000000000;
mem[757]  = 80'h00000000000000000000;
mem[758]  = 80'h00000000000000000000;
mem[759]  = 80'h10100000010000010010;
mem[760]  = 80'h00109400000208004500;
mem[761]  = 80'h0010002e292b0000fffd;
mem[762]  = 80'h0010104fc0550102c000;
mem[763]  = 80'h00100001ffabffabffab;
mem[764]  = 80'h0010d4d3f633d9ed3889;
mem[765]  = 80'h0010c8826f5ee365aa70;
mem[766]  = 80'h01104aef11da19f566ac;
mem[767]  = 80'h00000000000000000000;
mem[768]  = 80'h10100000010000010010;
mem[769]  = 80'h00109400000208004500;
mem[770]  = 80'h0010002e292c0000fffd;
mem[771]  = 80'h0010104ec0550102c000;
mem[772]  = 80'h00100001ffabffabffab;
mem[773]  = 80'h0010d3f732d908f9b709;
mem[774]  = 80'h0010706d7e32df84d895;
mem[775]  = 80'h0110618b30e628399323;
mem[776]  = 80'h00000000000000000000;
mem[777]  = 80'h00000000000000000000;
mem[778]  = 80'h00000000000000000000;
mem[779]  = 80'h00000000000000000000;
mem[780]  = 80'h10100000010000010010;
mem[781]  = 80'h00109400000208004500;
mem[782]  = 80'h0010002e292d0000fffd;
mem[783]  = 80'h0010104dc0550102c000;
mem[784]  = 80'h00100001ffabffabffab;
mem[785]  = 80'h0010d286ecf5d08075b6;
mem[786]  = 80'h0010bbbff9df2a54a6c4;
mem[787]  = 80'h01103b17387ccd2d9d3f;
mem[788]  = 80'h00000000000000000000;
mem[789]  = 80'h00000000000000000000;
mem[790]  = 80'h00000000000000000000;
mem[791]  = 80'h10100000010000010010;
mem[792]  = 80'h00109400000208004500;
mem[793]  = 80'h0010002e292e0000fffd;
mem[794]  = 80'h0010104cc0550102c000;
mem[795]  = 80'h00100001ffabffabffab;
mem[796]  = 80'h0010d1148e80b80a3276;
mem[797]  = 80'h0010e7c871e93424ef36;
mem[798]  = 80'h01100e3c2aa047965fb4;
mem[799]  = 80'h00000000000000000000;
mem[800]  = 80'h10100000010000010010;
mem[801]  = 80'h00109400000208004500;
mem[802]  = 80'h0010002e292f0000fffd;
mem[803]  = 80'h0010104bc0550102c000;
mem[804]  = 80'h00100001ffabffabffab;
mem[805]  = 80'h0010d06550ac6073f0c9;
mem[806]  = 80'h00102c1af604c1f4a667;
mem[807]  = 80'h0110c8a23a92e4dfb097;
mem[808]  = 80'h00000000000000000000;
mem[809]  = 80'h00000000000000000000;
mem[810]  = 80'h00000000000000000000;
mem[811]  = 80'h10100000010000010010;
mem[812]  = 80'h00109400000208004500;
mem[813]  = 80'h0010002e29300000fffd;
mem[814]  = 80'h0010104ac0550102c000;
mem[815]  = 80'h00100001ffabffabffab;
mem[816]  = 80'h0010cf6421724cab890b;
mem[817]  = 80'h001093d13b822c010c02;
mem[818]  = 80'h0110ef3542e54a4e60b7;
mem[819]  = 80'h00000000000000000000;
mem[820]  = 80'h00000000000000000000;
mem[821]  = 80'h00000000000000000000;
mem[822]  = 80'h10100000010000010010;
mem[823]  = 80'h00109400000208004500;
mem[824]  = 80'h0010002e29310000fffd;
mem[825]  = 80'h00101049c0550102c000;
mem[826]  = 80'h00100001ffabffabffab;
mem[827]  = 80'h0010ce15ff5e94d24bb4;
mem[828]  = 80'h00105803bc6fd9d14d53;
mem[829]  = 80'h0110a002766955368f6b;
mem[830]  = 80'h00000000000000000000;
mem[831]  = 80'h00000000000000000000;
mem[832]  = 80'h00000000000000000000;
mem[833]  = 80'h10100000010000010010;
mem[834]  = 80'h00109400000208004500;
mem[835]  = 80'h0010002e29320000fffd;
mem[836]  = 80'h00101048c0550102c000;
mem[837]  = 80'h00100001ffabffabffab;
mem[838]  = 80'h0010cd879d2bfc580c74;
mem[839]  = 80'h001004743459c7ae0ca1;
mem[840]  = 80'h011030b14eb11577e51b;
mem[841]  = 80'h00000000000000000000;
mem[842]  = 80'h10100000010000010010;
mem[843]  = 80'h00109400000208004500;
mem[844]  = 80'h0010002e29330000fffd;
mem[845]  = 80'h00101047c0550102c000;
mem[846]  = 80'h00100001ffabffabffab;
mem[847]  = 80'h0010ccf643072421cecb;
mem[848]  = 80'h0010cfa6b3b4327e4cf0;
mem[849]  = 80'h01104cb7ad93d72ba976;
mem[850]  = 80'h00000000000000000000;
mem[851]  = 80'h00000000000000000000;
mem[852]  = 80'h00000000000000000000;
mem[853]  = 80'h10100000010000010010;
mem[854]  = 80'h00109400000208004500;
mem[855]  = 80'h0010002e29340000fffd;
mem[856]  = 80'h00101046c0550102c000;
mem[857]  = 80'h00100001ffabffabffab;
mem[858]  = 80'h0010cbd287edf535414b;
mem[859]  = 80'h00107749a2d80e9f0815;
mem[860]  = 80'h0110c8e07c07ab9bebd4;
mem[861]  = 80'h00000000000000000000;
mem[862]  = 80'h00000000000000000000;
mem[863]  = 80'h00000000000000000000;
mem[864]  = 80'h10100000010000010010;
mem[865]  = 80'h00109400000208004500;
mem[866]  = 80'h0010002e29350000fffd;
mem[867]  = 80'h00101045c0550102c000;
mem[868]  = 80'h00100001ffabffabffab;
mem[869]  = 80'h0010caa359c12d4c83f4;
mem[870]  = 80'h0010bc9b2535fb4f0044;
mem[871]  = 80'h011030831c72b79af5d1;
mem[872]  = 80'h00000000000000000000;
mem[873]  = 80'h00000000000000000000;
mem[874]  = 80'h00000000000000000000;
mem[875]  = 80'h10100000010000010010;
mem[876]  = 80'h00109400000208004500;
mem[877]  = 80'h0010002e29360000fffd;
mem[878]  = 80'h00101044c0550102c000;
mem[879]  = 80'h00100001ffabffabffab;
mem[880]  = 80'h0010c9313bb445c6c434;
mem[881]  = 80'h0010e0ecad03e53f89b6;
mem[882]  = 80'h011013fce03b0f088015;
mem[883]  = 80'h00000000000000000000;
mem[884]  = 80'h10100000010000010010;
mem[885]  = 80'h00109400000208004500;
mem[886]  = 80'h0010002e29370000fffd;
mem[887]  = 80'h00101043c0550102c000;
mem[888]  = 80'h00100001ffabffabffab;
mem[889]  = 80'h0010c840e5989dbf068b;
mem[890]  = 80'h00102b3e2aee10ef10e7;
mem[891]  = 80'h0110c04575931fbcba28;
mem[892]  = 80'h00000000000000000000;
mem[893]  = 80'h00000000000000000000;
mem[894]  = 80'h00000000000000000000;
mem[895]  = 80'h00000000000000000000;
mem[896]  = 80'h10100000010000010010;
mem[897]  = 80'h00109400000208004500;
mem[898]  = 80'h0010002e29380000fffd;
mem[899]  = 80'h00101042c0550102c000;
mem[900]  = 80'h00100001ffabffabffab;
mem[901]  = 80'h0010c778b261e7efdb35;
mem[902]  = 80'h001091328fdb9cfdee7d;
mem[903]  = 80'h011028efed864c5c6ab2;
mem[904]  = 80'h00000000000000000000;
mem[905]  = 80'h00000000000000000000;
mem[906]  = 80'h00000000000000000000;
mem[907]  = 80'h10100000010000010010;
mem[908]  = 80'h00109400000208004500;
mem[909]  = 80'h0010002e29390000fffd;
mem[910]  = 80'h00101041c0550102c000;
mem[911]  = 80'h00100001ffabffabffab;
mem[912]  = 80'h0010c6096c4d3f96198a;
mem[913]  = 80'h00105ae00836692de12c;
mem[914]  = 80'h0110491b7dfc9f916616;
mem[915]  = 80'h00000000000000000000;
mem[916]  = 80'h10100000010000010010;
mem[917]  = 80'h00109400000208004500;
mem[918]  = 80'h0010002e293a0000fffd;
mem[919]  = 80'h00101040c0550102c000;
mem[920]  = 80'h00100001ffabffabffab;
mem[921]  = 80'h0010c59b0e38571c5e4a;
mem[922]  = 80'h001006978000775d52de;
mem[923]  = 80'h0110803aa5b78005f4b7;
mem[924]  = 80'h00000000000000000000;
mem[925]  = 80'h00000000000000000000;
mem[926]  = 80'h00000000000000000000;
mem[927]  = 80'h10100000010000010010;
mem[928]  = 80'h00109400000208004500;
mem[929]  = 80'h0010002e293b0000fffd;
mem[930]  = 80'h0010103fc0550102c000;
mem[931]  = 80'h00100001ffabffabffab;
mem[932]  = 80'h0010c4ead0148f659cf5;
mem[933]  = 80'h0010cd4507ed828d118f;
mem[934]  = 80'h0110a96f2be649aacce3;
mem[935]  = 80'h00000000000000000000;
mem[936]  = 80'h00000000000000000000;
mem[937]  = 80'h00000000000000000000;
mem[938]  = 80'h10100000010000010010;
mem[939]  = 80'h00109400000208004500;
mem[940]  = 80'h0010002e293c0000fffd;
mem[941]  = 80'h0010103ec0550102c000;
mem[942]  = 80'h00100001ffabffabffab;
mem[943]  = 80'h0010c3ce14fe5e711375;
mem[944]  = 80'h001075aa1681be6da26a;
mem[945]  = 80'h0110905e37ea80abaccc;
mem[946]  = 80'h00000000000000000000;
mem[947]  = 80'h00000000000000000000;
mem[948]  = 80'h00000000000000000000;
mem[949]  = 80'h10100000010000010010;
mem[950]  = 80'h00109400000208004500;
mem[951]  = 80'h0010002e293d0000fffd;
mem[952]  = 80'h0010103dc0550102c000;
mem[953]  = 80'h00100001ffabffabffab;
mem[954]  = 80'h0010c2bfcad28608d1ca;
mem[955]  = 80'h0010be78916c4bbdfd3b;
mem[956]  = 80'h0110ff1582a57eb4b3f4;
mem[957]  = 80'h00000000000000000000;
mem[958]  = 80'h10100000010000010010;
mem[959]  = 80'h00109400000208004500;
mem[960]  = 80'h0010002e293e0000fffd;
mem[961]  = 80'h0010103cc0550102c000;
mem[962]  = 80'h00100001ffabffabffab;
mem[963]  = 80'h0010c12da8a7ee82960a;
mem[964]  = 80'h0010e20f195a55cd35c9;
mem[965]  = 80'h0110e297a804cd989920;
mem[966]  = 80'h00000000000000000000;
mem[967]  = 80'h00000000000000000000;
mem[968]  = 80'h00000000000000000000;
mem[969]  = 80'h10100000010000010010;
mem[970]  = 80'h00109400000208004500;
mem[971]  = 80'h0010002e293f0000fffd;
mem[972]  = 80'h0010103bc0550102c000;
mem[973]  = 80'h00100001ffabffabffab;
mem[974]  = 80'h0010c05c768b36fb54b5;
mem[975]  = 80'h001029dd9eb7a01d7d98;
mem[976]  = 80'h011017383fe457670213;
mem[977]  = 80'h00000000000000000000;
mem[978]  = 80'h00000000000000000000;
mem[979]  = 80'h00000000000000000000;
mem[980]  = 80'h10100000010000010010;
mem[981]  = 80'h00109400000208004500;
mem[982]  = 80'h0010002e29400000fffd;
mem[983]  = 80'h0010103ac0550102c000;
mem[984]  = 80'h00100001ffabffabffab;
mem[985]  = 80'h0010bfcbd386ed10f47f;
mem[986]  = 80'h00108a85209a09ba88ff;
mem[987]  = 80'h011067d8e56a9079ae9f;
mem[988]  = 80'h00000000000000000000;
mem[989]  = 80'h00000000000000000000;
mem[990]  = 80'h00000000000000000000;
mem[991]  = 80'h10100000010000010010;
mem[992]  = 80'h00109400000208004500;
mem[993]  = 80'h0010002e29410000fffd;
mem[994]  = 80'h00101039c0550102c000;
mem[995]  = 80'h00100001ffabffabffab;
mem[996]  = 80'h0010beba0daa356936c0;
mem[997]  = 80'h00104157a777fc6a0bae;
mem[998]  = 80'h011058d97db0aa8002d4;
mem[999]  = 80'h00000000000000000000;
mem[1000] = 80'h10100000010000010010;
mem[1001] = 80'h00109400000208004500;
mem[1002] = 80'h0010002e29420000fffd;
mem[1003] = 80'h00101038c0550102c000;
mem[1004] = 80'h00100001ffabffabffab;
mem[1005] = 80'h0010bd286fdf5de37100;
mem[1006] = 80'h00101d202f41e21a885c;
mem[1007] = 80'h0110946db8cdb4603a8d;
mem[1008] = 80'h00000000000000000000;
mem[1009] = 80'h00000000000000000000;
mem[1010] = 80'h00000000000000000000;
mem[1011] = 80'h00000000000000000000;
mem[1012] = 80'h10100000010000010010;
mem[1013] = 80'h00109400000208004500;
mem[1014] = 80'h0010002e29430000fffd;
mem[1015] = 80'h00101037c0550102c000;
mem[1016] = 80'h00100001ffabffabffab;
mem[1017] = 80'h0010bc59b1f3859ab3bf;
mem[1018] = 80'h0010d6f2a8ac17ca890d;
mem[1019] = 80'h0110d696614ab0038f0a;
mem[1020] = 80'h00000000000000000000;
mem[1021] = 80'h00000000000000000000;
mem[1022] = 80'h00000000000000000000;
mem[1023] = 80'h10100000010000010010;
mem[1024] = 80'h00109400000208004500;
mem[1025] = 80'h0010002e29440000fffd;
mem[1026] = 80'h00101036c0550102c000;
mem[1027] = 80'h00100001ffabffabffab;
mem[1028] = 80'h0010bb7d7519548e3c3f;
mem[1029] = 80'h00106e1db9c02b2bece8;
mem[1030] = 80'h011067169792a7f1a18e;
mem[1031] = 80'h00000000000000000000;
mem[1032] = 80'h10100000010000010010;
mem[1033] = 80'h00109400000208004500;
mem[1034] = 80'h0010002e29450000fffd;
mem[1035] = 80'h00101035c0550102c000;
mem[1036] = 80'h00100001ffabffabffab;
mem[1037] = 80'h0010ba0cab358cf7fe80;
mem[1038] = 80'h0010a5cf3e2ddef865b9;
mem[1039] = 80'h0110ee8cf808db4100b1;
mem[1040] = 80'h00000000000000000000;
mem[1041] = 80'h00000000000000000000;
mem[1042] = 80'h00000000000000000000;
mem[1043] = 80'h10100000010000010010;
mem[1044] = 80'h00109400000208004500;
mem[1045] = 80'h0010002e29460000fffd;
mem[1046] = 80'h00101034c0550102c000;
mem[1047] = 80'h00100001ffabffabffab;
mem[1048] = 80'h0010b99ec940e47db940;
mem[1049] = 80'h0010f9b8b61bc088ec4b;
mem[1050] = 80'h0110cdf3b4c4740a620c;
mem[1051] = 80'h00000000000000000000;
mem[1052] = 80'h10100000010000010010;
mem[1053] = 80'h00109400000208004500;
mem[1054] = 80'h0010002e29470000fffd;
mem[1055] = 80'h00101033c0550102c000;
mem[1056] = 80'h00100001ffabffabffab;
mem[1057] = 80'h0010b8ef176c3c047bff;
mem[1058] = 80'h0010326a31f63558941a;
mem[1059] = 80'h01103dc90c04cf60f7de;
mem[1060] = 80'h00000000000000000000;
mem[1061] = 80'h00000000000000000000;
mem[1062] = 80'h00000000000000000000;
mem[1063] = 80'h00000000000000000000;
mem[1064] = 80'h10100000010000010010;
mem[1065] = 80'h00109400000208004500;
mem[1066] = 80'h0010002e29480000fffd;
mem[1067] = 80'h00101032c0550102c000;
mem[1068] = 80'h00100001ffabffabffab;
mem[1069] = 80'h0010b7d740954654a641;
mem[1070] = 80'h0010886694c3b94a2580;
mem[1071] = 80'h0110c8915676ee510084;
mem[1072] = 80'h00000000000000000000;
mem[1073] = 80'h00000000000000000000;
mem[1074] = 80'h00000000000000000000;
mem[1075] = 80'h10100000010000010010;
mem[1076] = 80'h00109400000208004500;
mem[1077] = 80'h0010002e29490000fffd;
mem[1078] = 80'h00101031c0550102c000;
mem[1079] = 80'h00100001ffabffabffab;
mem[1080] = 80'h0010b6a69eb99e2d64fe;
mem[1081] = 80'h001043b4132e4c9a65d1;
mem[1082] = 80'h0110b497e98da3879242;
mem[1083] = 80'h00000000000000000000;
mem[1084] = 80'h00000000000000000000;
mem[1085] = 80'h00000000000000000000;
mem[1086] = 80'h10100000010000010010;
mem[1087] = 80'h00109400000208004500;
mem[1088] = 80'h0010002e294a0000fffd;
mem[1089] = 80'h00101030c0550102c000;
mem[1090] = 80'h00100001ffabffabffab;
mem[1091] = 80'h0010b534fcccf6a7233e;
mem[1092] = 80'h00101fc39b1852ea3423;
mem[1093] = 80'h01100b66e6c89a1d9052;
mem[1094] = 80'h00000000000000000000;
mem[1095] = 80'h10100000010000010010;
mem[1096] = 80'h00109400000208004500;
mem[1097] = 80'h0010002e294b0000fffd;
mem[1098] = 80'h0010102fc0550102c000;
mem[1099] = 80'h00100001ffabffabffab;
mem[1100] = 80'h0010b44522e02edee181;
mem[1101] = 80'h0010d4111cf5a73a7572;
mem[1102] = 80'h01104451c67490342d8b;
mem[1103] = 80'h00000000000000000000;
mem[1104] = 80'h00000000000000000000;
mem[1105] = 80'h00000000000000000000;
mem[1106] = 80'h10100000010000010010;
mem[1107] = 80'h00109400000208004500;
mem[1108] = 80'h0010002e294c0000fffd;
mem[1109] = 80'h0010102ec0550102c000;
mem[1110] = 80'h00100001ffabffabffab;
mem[1111] = 80'h0010b361e60affca6e01;
mem[1112] = 80'h00106cfe0d999bdb4097;
mem[1113] = 80'h0110fb6ea64d1cff46dd;
mem[1114] = 80'h00000000000000000000;
mem[1115] = 80'h10100000010000010010;
mem[1116] = 80'h00109400000208004500;
mem[1117] = 80'h0010002e294d0000fffd;
mem[1118] = 80'h0010102dc0550102c000;
mem[1119] = 80'h00100001ffabffabffab;
mem[1120] = 80'h0010b210382627b3acbe;
mem[1121] = 80'h0010a72c8a746e0b39c6;
mem[1122] = 80'h011038652f7fca59cc1e;
mem[1123] = 80'h00000000000000000000;
mem[1124] = 80'h00000000000000000000;
mem[1125] = 80'h00000000000000000000;
mem[1126] = 80'h00000000000000000000;
mem[1127] = 80'h10100000010000010010;
mem[1128] = 80'h00109400000208004500;
mem[1129] = 80'h0010002e294e0000fffd;
mem[1130] = 80'h0010102cc0550102c000;
mem[1131] = 80'h00100001ffabffabffab;
mem[1132] = 80'h0010b1825a534f39eb7e;
mem[1133] = 80'h0010fb5b0242707bb034;
mem[1134] = 80'h01101b1a8009d8e849fd;
mem[1135] = 80'h00000000000000000000;
mem[1136] = 80'h00000000000000000000;
mem[1137] = 80'h00000000000000000000;
mem[1138] = 80'h00000000000000000000;
mem[1139] = 80'h10100000010000010010;
mem[1140] = 80'h00109400000208004500;
mem[1141] = 80'h0010002e294f0000fffd;
mem[1142] = 80'h0010102bc0550102c000;
mem[1143] = 80'h00100001ffabffabffab;
mem[1144] = 80'h0010b0f3847f974029c1;
mem[1145] = 80'h0010308985af85aa3965;
mem[1146] = 80'h0110fce09761f13196fa;
mem[1147] = 80'h00000000000000000000;
mem[1148] = 80'h00000000000000000000;
mem[1149] = 80'h00000000000000000000;
mem[1150] = 80'h10100000010000010010;
mem[1151] = 80'h00109400000208004500;
mem[1152] = 80'h0010002e29500000fffd;
mem[1153] = 80'h0010102ac0550102c000;
mem[1154] = 80'h00100001ffabffabffab;
mem[1155] = 80'h0010aff2f5a1bb985003;
mem[1156] = 80'h00108f424829685fcd00;
mem[1157] = 80'h0110f6c74b3bb36570f4;
mem[1158] = 80'h00000000000000000000;
mem[1159] = 80'h10100000010000010010;
mem[1160] = 80'h00109400000208004500;
mem[1161] = 80'h0010002e29510000fffd;
mem[1162] = 80'h00101029c0550102c000;
mem[1163] = 80'h00100001ffabffabffab;
mem[1164] = 80'h0010ae832b8d63e192bc;
mem[1165] = 80'h00104490cfc49d8fd251;
mem[1166] = 80'h0110944016dad330210e;
mem[1167] = 80'h00000000000000000000;
mem[1168] = 80'h00000000000000000000;
mem[1169] = 80'h00000000000000000000;
mem[1170] = 80'h10100000010000010010;
mem[1171] = 80'h00109400000208004500;
mem[1172] = 80'h0010002e29520000fffd;
mem[1173] = 80'h00101028c0550102c000;
mem[1174] = 80'h00100001ffabffabffab;
mem[1175] = 80'h0010ad1149f80b6bd57c;
mem[1176] = 80'h001018e747f283ff52a3;
mem[1177] = 80'h01100da7e2ea85f7948d;
mem[1178] = 80'h00000000000000000000;
mem[1179] = 80'h10100000010000010010;
mem[1180] = 80'h00109400000208004500;
mem[1181] = 80'h0010002e29530000fffd;
mem[1182] = 80'h00101027c0550102c000;
mem[1183] = 80'h00100001ffabffabffab;
mem[1184] = 80'h0010ac6097d4d31217c3;
mem[1185] = 80'h0010d335c01f762fd2f2;
mem[1186] = 80'h011067f58c87db81b987;
mem[1187] = 80'h00000000000000000000;
mem[1188] = 80'h00000000000000000000;
mem[1189] = 80'h00000000000000000000;
mem[1190] = 80'h10100000010000010010;
mem[1191] = 80'h00109400000208004500;
mem[1192] = 80'h0010002e29540000fffd;
mem[1193] = 80'h00101026c0550102c000;
mem[1194] = 80'h00100001ffabffabffab;
mem[1195] = 80'h0010ab44533e02069843;
mem[1196] = 80'h00106bdad1734ace9617;
mem[1197] = 80'h0110e3a2655c5dd107d4;
mem[1198] = 80'h00000000000000000000;
mem[1199] = 80'h00000000000000000000;
mem[1200] = 80'h00000000000000000000;
mem[1201] = 80'h10100000010000010010;
mem[1202] = 80'h00109400000208004500;
mem[1203] = 80'h0010002e29550000fffd;
mem[1204] = 80'h00101025c0550102c000;
mem[1205] = 80'h00100001ffabffabffab;
mem[1206] = 80'h0010aa358d12da7f5afc;
mem[1207] = 80'h0010a008569ebf1edd46;
mem[1208] = 80'h0110435ebcd04a2f4551;
mem[1209] = 80'h00000000000000000000;
mem[1210] = 80'h00000000000000000000;
mem[1211] = 80'h00000000000000000000;
mem[1212] = 80'h10100000010000010010;
mem[1213] = 80'h00109400000208004500;
mem[1214] = 80'h0010002e29560000fffd;
mem[1215] = 80'h00101024c0550102c000;
mem[1216] = 80'h00100001ffabffabffab;
mem[1217] = 80'h0010a9a7ef67b2f51d3c;
mem[1218] = 80'h0010fc7fdea8a16e16b4;
mem[1219] = 80'h01100b8ff7e3a0b635f3;
mem[1220] = 80'h00000000000000000000;
mem[1221] = 80'h10100000010000010010;
mem[1222] = 80'h00109400000208004500;
mem[1223] = 80'h0010002e29570000fffd;
mem[1224] = 80'h00101023c0550102c000;
mem[1225] = 80'h00100001ffabffabffab;
mem[1226] = 80'h0010a8d6314b6a8cdf83;
mem[1227] = 80'h001037ad594554be49e5;
mem[1228] = 80'h011064c44773fcc1ab28;
mem[1229] = 80'h00000000000000000000;
mem[1230] = 80'h00000000000000000000;
mem[1231] = 80'h00000000000000000000;
mem[1232] = 80'h00000000000000000000;
mem[1233] = 80'h10100000010000010010;
mem[1234] = 80'h00109400000208004500;
mem[1235] = 80'h0010002e29580000fffd;
mem[1236] = 80'h00101022c0550102c000;
mem[1237] = 80'h00100001ffabffabffab;
mem[1238] = 80'h0010a7ee66b210dc023d;
mem[1239] = 80'h00108da1fc70d8ab7f7f;
mem[1240] = 80'h011096036604f5797763;
mem[1241] = 80'h00000000000000000000;
mem[1242] = 80'h00000000000000000000;
mem[1243] = 80'h00000000000000000000;
mem[1244] = 80'h10100000010000010010;
mem[1245] = 80'h00109400000208004500;
mem[1246] = 80'h0010002e29590000fffd;
mem[1247] = 80'h00101021c0550102c000;
mem[1248] = 80'h00100001ffabffabffab;
mem[1249] = 80'h0010a69fb89ec8a5c082;
mem[1250] = 80'h001046737b9d2d7b3c2e;
mem[1251] = 80'h0110bf562c880843f216;
mem[1252] = 80'h00000000000000000000;
mem[1253] = 80'h10100000010000010010;
mem[1254] = 80'h00109400000208004500;
mem[1255] = 80'h0010002e295a0000fffd;
mem[1256] = 80'h00101020c0550102c000;
mem[1257] = 80'h00100001ffabffabffab;
mem[1258] = 80'h0010a50ddaeba02f8742;
mem[1259] = 80'h00101a04f3ab330b8fdc;
mem[1260] = 80'h0110767711851b34d60b;
mem[1261] = 80'h00000000000000000000;
mem[1262] = 80'h00000000000000000000;
mem[1263] = 80'h00000000000000000000;
mem[1264] = 80'h00000000000000000000;
mem[1265] = 80'h10100000010000010010;
mem[1266] = 80'h00109400000208004500;
mem[1267] = 80'h0010002e295b0000fffd;
mem[1268] = 80'h0010101fc0550102c000;
mem[1269] = 80'h00100001ffabffabffab;
mem[1270] = 80'h0010a47c04c7785645fd;
mem[1271] = 80'h0010d1d67446c6db8e8d;
mem[1272] = 80'h0110348cc855955f62a9;
mem[1273] = 80'h00000000000000000000;
mem[1274] = 80'h00000000000000000000;
mem[1275] = 80'h00000000000000000000;
mem[1276] = 80'h10100000010000010010;
mem[1277] = 80'h00109400000208004500;
mem[1278] = 80'h0010002e295c0000fffd;
mem[1279] = 80'h0010101ec0550102c000;
mem[1280] = 80'h00100001ffabffabffab;
mem[1281] = 80'h0010a358c02da942ca7d;
mem[1282] = 80'h00106939652afa3afb68;
mem[1283] = 80'h0110867fde31b5da31f6;
mem[1284] = 80'h00000000000000000000;
mem[1285] = 80'h10100000010000010010;
mem[1286] = 80'h00109400000208004500;
mem[1287] = 80'h0010002e295d0000fffd;
mem[1288] = 80'h0010101dc0550102c000;
mem[1289] = 80'h00100001ffabffabffab;
mem[1290] = 80'h0010a2291e01713b08c2;
mem[1291] = 80'h0010a2ebe2c70fea6339;
mem[1292] = 80'h011066f76609e1ffdf9f;
mem[1293] = 80'h00000000000000000000;
mem[1294] = 80'h00000000000000000000;
mem[1295] = 80'h00000000000000000000;
mem[1296] = 80'h10100000010000010010;
mem[1297] = 80'h00109400000208004500;
mem[1298] = 80'h0010002e295e0000fffd;
mem[1299] = 80'h0010101cc0550102c000;
mem[1300] = 80'h00100001ffabffabffab;
mem[1301] = 80'h0010a1bb7c7419b14f02;
mem[1302] = 80'h0010fe9c6af1119aebcb;
mem[1303] = 80'h011076b99b6e9a5a0c92;
mem[1304] = 80'h00000000000000000000;
mem[1305] = 80'h00000000000000000000;
mem[1306] = 80'h00000000000000000000;
mem[1307] = 80'h10100000010000010010;
mem[1308] = 80'h00109400000208004500;
mem[1309] = 80'h0010002e295f0000fffd;
mem[1310] = 80'h0010101bc0550102c000;
mem[1311] = 80'h00100001ffabffabffab;
mem[1312] = 80'h0010a0caa258c1c88dbd;
mem[1313] = 80'h0010354eed1ce44ae39a;
mem[1314] = 80'h01108edaf42ad114cec9;
mem[1315] = 80'h00000000000000000000;
mem[1316] = 80'h00000000000000000000;
mem[1317] = 80'h00000000000000000000;
mem[1318] = 80'h10100000010000010010;
mem[1319] = 80'h00109400000208004500;
mem[1320] = 80'h0010002e29600000fffd;
mem[1321] = 80'h0010101ac0550102c000;
mem[1322] = 80'h00100001ffabffabffab;
mem[1323] = 80'h00109fb99fc84001bc87;
mem[1324] = 80'h0010810bf1fcca713c01;
mem[1325] = 80'h0110775cd31c3722d895;
mem[1326] = 80'h00000000000000000000;
mem[1327] = 80'h10100000010000010010;
mem[1328] = 80'h00109400000208004500;
mem[1329] = 80'h0010002e29610000fffd;
mem[1330] = 80'h00101019c0550102c000;
mem[1331] = 80'h00100001ffabffabffab;
mem[1332] = 80'h00109ec841e498787e38;
mem[1333] = 80'h00104ad976113fa17d50;
mem[1334] = 80'h0110386b525a7b2b34ab;
mem[1335] = 80'h00000000000000000000;
mem[1336] = 80'h00000000000000000000;
mem[1337] = 80'h00000000000000000000;
mem[1338] = 80'h10100000010000010010;
mem[1339] = 80'h00109400000208004500;
mem[1340] = 80'h0010002e29620000fffd;
mem[1341] = 80'h00101018c0550102c000;
mem[1342] = 80'h00100001ffabffabffab;
mem[1343] = 80'h00109d5a2391f0f239f8;
mem[1344] = 80'h001016aefe2721d03ca2;
mem[1345] = 80'h0110b3d9ed067ae2ac93;
mem[1346] = 80'h00000000000000000000;
mem[1347] = 80'h00000000000000000000;
mem[1348] = 80'h00000000000000000000;
mem[1349] = 80'h10100000010000010010;
mem[1350] = 80'h00109400000208004500;
mem[1351] = 80'h0010002e29630000fffd;
mem[1352] = 80'h00101017c0550102c000;
mem[1353] = 80'h00100001ffabffabffab;
mem[1354] = 80'h00109c2bfdbd288bfb47;
mem[1355] = 80'h0010dd7c79cad4007df3;
mem[1356] = 80'h0110fcee9c18ea21939e;
mem[1357] = 80'h00000000000000000000;
mem[1358] = 80'h00000000000000000000;
mem[1359] = 80'h00000000000000000000;
mem[1360] = 80'h10100000010000010010;
mem[1361] = 80'h00109400000208004500;
mem[1362] = 80'h0010002e29640000fffd;
mem[1363] = 80'h00101016c0550102c000;
mem[1364] = 80'h00100001ffabffabffab;
mem[1365] = 80'h00109b0f3957f99f74c7;
mem[1366] = 80'h0010659368a6e8e15816;
mem[1367] = 80'h011040a26d5d5617c5be;
mem[1368] = 80'h00000000000000000000;
mem[1369] = 80'h10100000010000010010;
mem[1370] = 80'h00109400000208004500;
mem[1371] = 80'h0010002e29650000fffd;
mem[1372] = 80'h00101015c0550102c000;
mem[1373] = 80'h00100001ffabffabffab;
mem[1374] = 80'h00109a7ee77b21e6b678;
mem[1375] = 80'h0010ae41ef4b1d311247;
mem[1376] = 80'h0110d36f05318d9f386a;
mem[1377] = 80'h00000000000000000000;
mem[1378] = 80'h00000000000000000000;
mem[1379] = 80'h00000000000000000000;
mem[1380] = 80'h00000000000000000000;
mem[1381] = 80'h10100000010000010010;
mem[1382] = 80'h00109400000208004500;
mem[1383] = 80'h0010002e29660000fffd;
mem[1384] = 80'h00101014c0550102c000;
mem[1385] = 80'h00100001ffabffabffab;
mem[1386] = 80'h001099ec850e496cf1b8;
mem[1387] = 80'h0010f236677d03415ab5;
mem[1388] = 80'h0110d57518bf5d036cef;
mem[1389] = 80'h00000000000000000000;
mem[1390] = 80'h10100000010000010010;
mem[1391] = 80'h00109400000208004500;
mem[1392] = 80'h0010002e29670000fffd;
mem[1393] = 80'h00101013c0550102c000;
mem[1394] = 80'h00100001ffabffabffab;
mem[1395] = 80'h0010989d5b2291153307;
mem[1396] = 80'h001039e4e090f69121e4;
mem[1397] = 80'h0110701ca51b3525ec1e;
mem[1398] = 80'h00000000000000000000;
mem[1399] = 80'h00000000000000000000;
mem[1400] = 80'h00000000000000000000;
mem[1401] = 80'h10100000010000010010;
mem[1402] = 80'h00109400000208004500;
mem[1403] = 80'h0010002e29680000fffd;
mem[1404] = 80'h00101012c0550102c000;
mem[1405] = 80'h00100001ffabffabffab;
mem[1406] = 80'h001097a50cdbeb45eeb9;
mem[1407] = 80'h001083e845a57a83d07e;
mem[1408] = 80'h01108888e4668a7f1518;
mem[1409] = 80'h00000000000000000000;
mem[1410] = 80'h00000000000000000000;
mem[1411] = 80'h00000000000000000000;
mem[1412] = 80'h10100000010000010010;
mem[1413] = 80'h00109400000208004500;
mem[1414] = 80'h0010002e29690000fffd;
mem[1415] = 80'h00101011c0550102c000;
mem[1416] = 80'h00100001ffabffabffab;
mem[1417] = 80'h001096d4d2f7333c2c06;
mem[1418] = 80'h0010483ac2488f53d02f;
mem[1419] = 80'h0110f942d3a7a3df568e;
mem[1420] = 80'h00000000000000000000;
mem[1421] = 80'h00000000000000000000;
mem[1422] = 80'h00000000000000000000;
mem[1423] = 80'h10100000010000010010;
mem[1424] = 80'h00109400000208004500;
mem[1425] = 80'h0010002e296a0000fffd;
mem[1426] = 80'h00101010c0550102c000;
mem[1427] = 80'h00100001ffabffabffab;
mem[1428] = 80'h00109546b0825bb66bc6;
mem[1429] = 80'h0010144d4a7e912340dd;
mem[1430] = 80'h011063d65e1716227259;
mem[1431] = 80'h00000000000000000000;
mem[1432] = 80'h00000000000000000000;
mem[1433] = 80'h00000000000000000000;
mem[1434] = 80'h10100000010000010010;
mem[1435] = 80'h00109400000208004500;
mem[1436] = 80'h0010002e296b0000fffd;
mem[1437] = 80'h0010100fc0550102c000;
mem[1438] = 80'h00100001ffabffabffab;
mem[1439] = 80'h001094376eae83cfa979;
mem[1440] = 80'h0010df9fcd9364f0cf8c;
mem[1441] = 80'h011040eaad3580e1c25a;
mem[1442] = 80'h00000000000000000000;
mem[1443] = 80'h10100000010000010010;
mem[1444] = 80'h00109400000208004500;
mem[1445] = 80'h0010002e296c0000fffd;
mem[1446] = 80'h0010100ec0550102c000;
mem[1447] = 80'h00100001ffabffabffab;
mem[1448] = 80'h00109313aa4452db26f9;
mem[1449] = 80'h00106770dcff5811b469;
mem[1450] = 80'h0110d11626d14a3517af;
mem[1451] = 80'h00000000000000000000;
mem[1452] = 80'h00000000000000000000;
mem[1453] = 80'h00000000000000000000;
mem[1454] = 80'h10100000010000010010;
mem[1455] = 80'h00109400000208004500;
mem[1456] = 80'h0010002e296d0000fffd;
mem[1457] = 80'h0010100dc0550102c000;
mem[1458] = 80'h00100001ffabffabffab;
mem[1459] = 80'h0010926274688aa2e446;
mem[1460] = 80'h0010aca25b12adc1cf38;
mem[1461] = 80'h0110747f911cf6718c18;
mem[1462] = 80'h00000000000000000000;
mem[1463] = 80'h00000000000000000000;
mem[1464] = 80'h00000000000000000000;
mem[1465] = 80'h10100000010000010010;
mem[1466] = 80'h00109400000208004500;
mem[1467] = 80'h0010002e296e0000fffd;
mem[1468] = 80'h0010100cc0550102c000;
mem[1469] = 80'h00100001ffabffabffab;
mem[1470] = 80'h001091f0161de228a386;
mem[1471] = 80'h0010f0d5d324b3b104ca;
mem[1472] = 80'h01103cae191eab6cf50b;
mem[1473] = 80'h00000000000000000000;
mem[1474] = 80'h10100000010000010010;
mem[1475] = 80'h00109400000208004500;
mem[1476] = 80'h0010002e296f0000fffd;
mem[1477] = 80'h0010100bc0550102c000;
mem[1478] = 80'h00100001ffabffabffab;
mem[1479] = 80'h00109081c8313a516139;
mem[1480] = 80'h00103b0754c946614b9b;
mem[1481] = 80'h01105096995eac842ace;
mem[1482] = 80'h00000000000000000000;
mem[1483] = 80'h00000000000000000000;
mem[1484] = 80'h00000000000000000000;
mem[1485] = 80'h10100000010000010010;
mem[1486] = 80'h00109400000208004500;
mem[1487] = 80'h0010002e29700000fffd;
mem[1488] = 80'h0010100ac0550102c000;
mem[1489] = 80'h00100001ffabffabffab;
mem[1490] = 80'h00108f80b9ef168918fb;
mem[1491] = 80'h001084cc994fab9466fe;
mem[1492] = 80'h0110f50e614de5351fd0;
mem[1493] = 80'h00000000000000000000;
mem[1494] = 80'h00000000000000000000;
mem[1495] = 80'h00000000000000000000;
mem[1496] = 80'h10100000010000010010;
mem[1497] = 80'h00109400000208004500;
mem[1498] = 80'h0010002e29710000fffd;
mem[1499] = 80'h00101009c0550102c000;
mem[1500] = 80'h00100001ffabffabffab;
mem[1501] = 80'h00108ef167c3cef0da44;
mem[1502] = 80'h00104f1e1ea25e4424af;
mem[1503] = 80'h0110ef6a7ff60a399bcf;
mem[1504] = 80'h00000000000000000000;
mem[1505] = 80'h00000000000000000000;
mem[1506] = 80'h00000000000000000000;
mem[1507] = 80'h10100000010000010010;
mem[1508] = 80'h00109400000208004500;
mem[1509] = 80'h0010002e29720000fffd;
mem[1510] = 80'h00101008c0550102c000;
mem[1511] = 80'h00100001ffabffabffab;
mem[1512] = 80'h00108d6305b6a67a9d84;
mem[1513] = 80'h0010136996944034e75d;
mem[1514] = 80'h01102e122945ef5294d5;
mem[1515] = 80'h00000000000000000000;
mem[1516] = 80'h00000000000000000000;
mem[1517] = 80'h00000000000000000000;
mem[1518] = 80'h10100000010000010010;
mem[1519] = 80'h00109400000208004500;
mem[1520] = 80'h0010002e29730000fffd;
mem[1521] = 80'h00101007c0550102c000;
mem[1522] = 80'h00100001ffabffabffab;
mem[1523] = 80'h00108c12db9a7e035f3b;
mem[1524] = 80'h0010d8bb1179b5e4a70c;
mem[1525] = 80'h0110521421d981ba8b29;
mem[1526] = 80'h00000000000000000000;
mem[1527] = 80'h10100000010000010010;
mem[1528] = 80'h00109400000208004500;
mem[1529] = 80'h0010002e29740000fffd;
mem[1530] = 80'h00101006c0550102c000;
mem[1531] = 80'h00100001ffabffabffab;
mem[1532] = 80'h00108b361f70af17d0bb;
mem[1533] = 80'h0010605400158905e3e9;
mem[1534] = 80'h0110d64331e9038b9388;
mem[1535] = 80'h00000000000000000000;
mem[1536] = 80'h00000000000000000000;
mem[1537] = 80'h00000000000000000000;
mem[1538] = 80'h10100000010000010010;
mem[1539] = 80'h00109400000208004500;
mem[1540] = 80'h0010002e29750000fffd;
mem[1541] = 80'h00101005c0550102c000;
mem[1542] = 80'h00100001ffabffabffab;
mem[1543] = 80'h00108a47c15c776e1204;
mem[1544] = 80'h0010ab8687f87cd46bb8;
mem[1545] = 80'h011002880c5520d068e5;
mem[1546] = 80'h00000000000000000000;
mem[1547] = 80'h00000000000000000000;
mem[1548] = 80'h00000000000000000000;
mem[1549] = 80'h10100000010000010010;
mem[1550] = 80'h00109400000208004500;
mem[1551] = 80'h0010002e29760000fffd;
mem[1552] = 80'h00101004c0550102c000;
mem[1553] = 80'h00100001ffabffabffab;
mem[1554] = 80'h001089d5a3291fe455c4;
mem[1555] = 80'h0010f7f10fce62a4e24a;
mem[1556] = 80'h011021f7eeb112a23b5d;
mem[1557] = 80'h00000000000000000000;
mem[1558] = 80'h00000000000000000000;
mem[1559] = 80'h00000000000000000000;
mem[1560] = 80'h10100000010000010010;
mem[1561] = 80'h00109400000208004500;
mem[1562] = 80'h0010002e29770000fffd;
mem[1563] = 80'h00101003c0550102c000;
mem[1564] = 80'h00100001ffabffabffab;
mem[1565] = 80'h001088a47d05c79d977b;
mem[1566] = 80'h00103c2388239774fb1b;
mem[1567] = 80'h0110e9d65a8e08285de8;
mem[1568] = 80'h00000000000000000000;
mem[1569] = 80'h10100000010000010010;
mem[1570] = 80'h00109400000208004500;
mem[1571] = 80'h0010002e29780000fffd;
mem[1572] = 80'h00101002c0550102c000;
mem[1573] = 80'h00100001ffabffabffab;
mem[1574] = 80'h0010879c2afcbdcd4ac5;
mem[1575] = 80'h0010862f2d161b660b81;
mem[1576] = 80'h0110227348347e205976;
mem[1577] = 80'h00000000000000000000;
mem[1578] = 80'h00000000000000000000;
mem[1579] = 80'h00000000000000000000;
mem[1580] = 80'h00000000000000000000;
mem[1581] = 80'h10100000010000010010;
mem[1582] = 80'h00109400000208004500;
mem[1583] = 80'h0010002e29790000fffd;
mem[1584] = 80'h00101001c0550102c000;
mem[1585] = 80'h00100001ffabffabffab;
mem[1586] = 80'h001086edf4d065b4887a;
mem[1587] = 80'h00104dfdaafbeeb68ad0;
mem[1588] = 80'h01107b10a881e940c81f;
mem[1589] = 80'h00000000000000000000;
mem[1590] = 80'h10100000010000010010;
mem[1591] = 80'h00109400000208004500;
mem[1592] = 80'h0010002e297a0000fffd;
mem[1593] = 80'h00101000c0550102c000;
mem[1594] = 80'h00100001ffabffabffab;
mem[1595] = 80'h0010857f96a50d3ecfba;
mem[1596] = 80'h0010118a22cdf0c63b22;
mem[1597] = 80'h0110d453d24d840a6149;
mem[1598] = 80'h00000000000000000000;
mem[1599] = 80'h00000000000000000000;
mem[1600] = 80'h00000000000000000000;
mem[1601] = 80'h10100000010000010010;
mem[1602] = 80'h00109400000208004500;
mem[1603] = 80'h0010002e297b0000fffd;
mem[1604] = 80'h00100fffc0550102c000;
mem[1605] = 80'h00100001ffabffabffab;
mem[1606] = 80'h0010840e4889d5470d05;
mem[1607] = 80'h0010da58a52005167573;
mem[1608] = 80'h01108b5acbbd24c9f4ca;
mem[1609] = 80'h00000000000000000000;
mem[1610] = 80'h00000000000000000000;
mem[1611] = 80'h00000000000000000000;
mem[1612] = 80'h10100000010000010010;
mem[1613] = 80'h00109400000208004500;
mem[1614] = 80'h0010002e297c0000fffd;
mem[1615] = 80'h00100ffec0550102c000;
mem[1616] = 80'h00100001ffabffabffab;
mem[1617] = 80'h0010832a8c6304538285;
mem[1618] = 80'h001062b7b44c39f74f96;
mem[1619] = 80'h0110245ba4ac4d9b08a1;
mem[1620] = 80'h00000000000000000000;
mem[1621] = 80'h00000000000000000000;
mem[1622] = 80'h00000000000000000000;
mem[1623] = 80'h10100000010000010010;
mem[1624] = 80'h00109400000208004500;
mem[1625] = 80'h0010002e297d0000fffd;
mem[1626] = 80'h00100ffdc0550102c000;
mem[1627] = 80'h00100001ffabffabffab;
mem[1628] = 80'h0010825b524fdc2a403a;
mem[1629] = 80'h0010a96533a1cc2715c7;
mem[1630] = 80'h0110b4e59b14b4b56546;
mem[1631] = 80'h00000000000000000000;
mem[1632] = 80'h00000000000000000000;
mem[1633] = 80'h00000000000000000000;
mem[1634] = 80'h10100000010000010010;
mem[1635] = 80'h00109400000208004500;
mem[1636] = 80'h0010002e297e0000fffd;
mem[1637] = 80'h00100ffcc0550102c000;
mem[1638] = 80'h00100001ffabffabffab;
mem[1639] = 80'h001081c9303ab4a007fa;
mem[1640] = 80'h0010f512bb97d2485e35;
mem[1641] = 80'h011088fe273a5febad2b;
mem[1642] = 80'h00000000000000000000;
mem[1643] = 80'h10100000010000010010;
mem[1644] = 80'h00109400000208004500;
mem[1645] = 80'h0010002e297f0000fffd;
mem[1646] = 80'h00100ffbc0550102c000;
mem[1647] = 80'h00100001ffabffabffab;
mem[1648] = 80'h001080b8ee166cd9c545;
mem[1649] = 80'h00103ec03c7a27981664;
mem[1650] = 80'h01107d5128899914cc53;
mem[1651] = 80'h00000000000000000000;
mem[1652] = 80'h00000000000000000000;
mem[1653] = 80'h00000000000000000000;
mem[1654] = 80'h00000000000000000000;
mem[1655] = 80'h10100000010000010010;
mem[1656] = 80'h00109400000208004500;
mem[1657] = 80'h0010002e29800000fffd;
mem[1658] = 80'h00100ffac0550102c000;
mem[1659] = 80'h00100001ffabffabffab;
mem[1660] = 80'h00107f97a40ddb0e84d0;
mem[1661] = 80'h00107871412174d7d1ab;
mem[1662] = 80'h0110b9aac2ba4f81a62f;
mem[1663] = 80'h00000000000000000000;
mem[1664] = 80'h10100000010000010010;
mem[1665] = 80'h00109400000208004500;
mem[1666] = 80'h0010002e29810000fffd;
mem[1667] = 80'h00100ff9c0550102c000;
mem[1668] = 80'h00100001ffabffabffab;
mem[1669] = 80'h00107ee67a210377466f;
mem[1670] = 80'h0010b3a3c6cc8107d2fa;
mem[1671] = 80'h01109d33516b3855847a;
mem[1672] = 80'h00000000000000000000;
mem[1673] = 80'h00000000000000000000;
mem[1674] = 80'h00000000000000000000;
mem[1675] = 80'h10100000010000010010;
mem[1676] = 80'h00109400000208004500;
mem[1677] = 80'h0010002e29820000fffd;
mem[1678] = 80'h00100ff8c0550102c000;
mem[1679] = 80'h00100001ffabffabffab;
mem[1680] = 80'h00107d7418546bfd01af;
mem[1681] = 80'h0010efd44efa9f775108;
mem[1682] = 80'h011051877bb4c19882c2;
mem[1683] = 80'h00000000000000000000;
mem[1684] = 80'h00000000000000000000;
mem[1685] = 80'h00000000000000000000;
mem[1686] = 80'h10100000010000010010;
mem[1687] = 80'h00109400000208004500;
mem[1688] = 80'h0010002e29830000fffd;
mem[1689] = 80'h00100ff7c0550102c000;
mem[1690] = 80'h00100001ffabffabffab;
mem[1691] = 80'h00107c05c678b384c310;
mem[1692] = 80'h00102406c9176aa7ce59;
mem[1693] = 80'h01102898f83457abaa35;
mem[1694] = 80'h00000000000000000000;
mem[1695] = 80'h00000000000000000000;
mem[1696] = 80'h00000000000000000000;
mem[1697] = 80'h10100000010000010010;
mem[1698] = 80'h00109400000208004500;
mem[1699] = 80'h0010002e29840000fffd;
mem[1700] = 80'h00100ff6c0550102c000;
mem[1701] = 80'h00100001ffabffabffab;
mem[1702] = 80'h00107b21029262904c90;
mem[1703] = 80'h00109ce9d87b5646b5bc;
mem[1704] = 80'h0110b964985e9dfbf577;
mem[1705] = 80'h00000000000000000000;
mem[1706] = 80'h10100000010000010010;
mem[1707] = 80'h00109400000208004500;
mem[1708] = 80'h0010002e29850000fffd;
mem[1709] = 80'h00100ff5c0550102c000;
mem[1710] = 80'h00100001ffabffabffab;
mem[1711] = 80'h00107a50dcbebae98e2f;
mem[1712] = 80'h0010573b5f96a396beed;
mem[1713] = 80'h01101454322da77d20be;
mem[1714] = 80'h00000000000000000000;
mem[1715] = 80'h00000000000000000000;
mem[1716] = 80'h00000000000000000000;
mem[1717] = 80'h00000000000000000000;
mem[1718] = 80'h10100000010000010010;
mem[1719] = 80'h00109400000208004500;
mem[1720] = 80'h0010002e29860000fffd;
mem[1721] = 80'h00100ff4c0550102c000;
mem[1722] = 80'h00100001ffabffabffab;
mem[1723] = 80'h001079c2becbd263c9ef;
mem[1724] = 80'h00100b4cd7a0bde6341f;
mem[1725] = 80'h01106278f3b297cdb06b;
mem[1726] = 80'h00000000000000000000;
mem[1727] = 80'h00000000000000000000;
mem[1728] = 80'h00000000000000000000;
mem[1729] = 80'h10100000010000010010;
mem[1730] = 80'h00109400000208004500;
mem[1731] = 80'h0010002e29870000fffd;
mem[1732] = 80'h00100ff3c0550102c000;
mem[1733] = 80'h00100001ffabffabffab;
mem[1734] = 80'h001078b360e70a1a0b50;
mem[1735] = 80'h0010c09e504d48364a4e;
mem[1736] = 80'h011038e434a676ef46b9;
mem[1737] = 80'h00000000000000000000;
mem[1738] = 80'h10100000010000010010;
mem[1739] = 80'h00109400000208004500;
mem[1740] = 80'h0010002e29880000fffd;
mem[1741] = 80'h00100ff2c0550102c000;
mem[1742] = 80'h00100001ffabffabffab;
mem[1743] = 80'h0010778b371e704ad6ee;
mem[1744] = 80'h00107a92f578c4257dd4;
mem[1745] = 80'h01104bb20c65f46c2ea4;
mem[1746] = 80'h00000000000000000000;
mem[1747] = 80'h00000000000000000000;
mem[1748] = 80'h00000000000000000000;
mem[1749] = 80'h10100000010000010010;
mem[1750] = 80'h00109400000208004500;
mem[1751] = 80'h0010002e29890000fffd;
mem[1752] = 80'h00100ff1c0550102c000;
mem[1753] = 80'h00100001ffabffabffab;
mem[1754] = 80'h001076fae932a8331451;
mem[1755] = 80'h0010b140729531f53e85;
mem[1756] = 80'h011062e7ec155dbc4831;
mem[1757] = 80'h00000000000000000000;
mem[1758] = 80'h00000000000000000000;
mem[1759] = 80'h00000000000000000000;
mem[1760] = 80'h00000000000000000000;
mem[1761] = 80'h10100000010000010010;
mem[1762] = 80'h00109400000208004500;
mem[1763] = 80'h0010002e298a0000fffd;
mem[1764] = 80'h00100ff0c0550102c000;
mem[1765] = 80'h00100001ffabffabffab;
mem[1766] = 80'h001075688b47c0b95391;
mem[1767] = 80'h0010ed37faa32f85ed77;
mem[1768] = 80'h0110a0ec453f567a6476;
mem[1769] = 80'h00000000000000000000;
mem[1770] = 80'h10100000010000010010;
mem[1771] = 80'h00109400000208004500;
mem[1772] = 80'h0010002e298b0000fffd;
mem[1773] = 80'h00100fefc0550102c000;
mem[1774] = 80'h00100001ffabffabffab;
mem[1775] = 80'h00107419556b18c0912e;
mem[1776] = 80'h001026e57d4eda55ac26;
mem[1777] = 80'h0110efdb72005005ebde;
mem[1778] = 80'h00000000000000000000;
mem[1779] = 80'h00000000000000000000;
mem[1780] = 80'h00000000000000000000;
mem[1781] = 80'h10100000010000010010;
mem[1782] = 80'h00109400000208004500;
mem[1783] = 80'h0010002e298c0000fffd;
mem[1784] = 80'h00100feec0550102c000;
mem[1785] = 80'h00100001ffabffabffab;
mem[1786] = 80'h0010733d9181c9d41eae;
mem[1787] = 80'h00109e0a6c22e6b419c3;
mem[1788] = 80'h01104b7cbc9cd2251074;
mem[1789] = 80'h00000000000000000000;
mem[1790] = 80'h00000000000000000000;
mem[1791] = 80'h00000000000000000000;
mem[1792] = 80'h10100000010000010010;
mem[1793] = 80'h00109400000208004500;
mem[1794] = 80'h0010002e298d0000fffd;
mem[1795] = 80'h00100fedc0550102c000;
mem[1796] = 80'h00100001ffabffabffab;
mem[1797] = 80'h0010724c4fad11addc11;
mem[1798] = 80'h001055d8ebcf13646092;
mem[1799] = 80'h011088771231b4bfef0d;
mem[1800] = 80'h00000000000000000000;
mem[1801] = 80'h00000000000000000000;
mem[1802] = 80'h00000000000000000000;
mem[1803] = 80'h10100000010000010010;
mem[1804] = 80'h00109400000208004500;
mem[1805] = 80'h0010002e298e0000fffd;
mem[1806] = 80'h00100fecc0550102c000;
mem[1807] = 80'h00100001ffabffabffab;
mem[1808] = 80'h001071de2dd879279bd1;
mem[1809] = 80'h001009af63f90d14e960;
mem[1810] = 80'h0110ab083c2a49baf1ff;
mem[1811] = 80'h00000000000000000000;
mem[1812] = 80'h10100000010000010010;
mem[1813] = 80'h00109400000208004500;
mem[1814] = 80'h0010002e298f0000fffd;
mem[1815] = 80'h00100febc0550102c000;
mem[1816] = 80'h00100001ffabffabffab;
mem[1817] = 80'h001070aff3f4a15e596e;
mem[1818] = 80'h0010c27de414f8c4e031;
mem[1819] = 80'h0110605ac0aa3f203d6e;
mem[1820] = 80'h00000000000000000000;
mem[1821] = 80'h00000000000000000000;
mem[1822] = 80'h00000000000000000000;
mem[1823] = 80'h10100000010000010010;
mem[1824] = 80'h00109400000208004500;
mem[1825] = 80'h0010002e29900000fffd;
mem[1826] = 80'h00100feac0550102c000;
mem[1827] = 80'h00100001ffabffabffab;
mem[1828] = 80'h00106fae822a8d8620ac;
mem[1829] = 80'h00107db6299215310a54;
mem[1830] = 80'h01104a014f255001f1c3;
mem[1831] = 80'h00000000000000000000;
mem[1832] = 80'h00000000000000000000;
mem[1833] = 80'h00000000000000000000;
mem[1834] = 80'h10100000010000010010;
mem[1835] = 80'h00109400000208004500;
mem[1836] = 80'h0010002e29910000fffd;
mem[1837] = 80'h00100fe9c0550102c000;
mem[1838] = 80'h00100001ffabffabffab;
mem[1839] = 80'h00106edf5c0655ffe213;
mem[1840] = 80'h0010b664ae7fe0e28805;
mem[1841] = 80'h01101f610fd9c84d8bf4;
mem[1842] = 80'h00000000000000000000;
mem[1843] = 80'h00000000000000000000;
mem[1844] = 80'h00000000000000000000;
mem[1845] = 80'h10100000010000010010;
mem[1846] = 80'h00109400000208004500;
mem[1847] = 80'h0010002e29920000fffd;
mem[1848] = 80'h00100fe8c0550102c000;
mem[1849] = 80'h00100001ffabffabffab;
mem[1850] = 80'h00106d4d3e733d75a5d3;
mem[1851] = 80'h0010ea132649fe920af7;
mem[1852] = 80'h0110e0e4762a08e9a8e3;
mem[1853] = 80'h00000000000000000000;
mem[1854] = 80'h10100000010000010010;
mem[1855] = 80'h00109400000208004500;
mem[1856] = 80'h0010002e29930000fffd;
mem[1857] = 80'h00100fe7c0550102c000;
mem[1858] = 80'h00100001ffabffabffab;
mem[1859] = 80'h00106c3ce05fe50c676c;
mem[1860] = 80'h001021c1a1a40b4274a6;
mem[1861] = 80'h0110ba7869232249fcd1;
mem[1862] = 80'h00000000000000000000;
mem[1863] = 80'h00000000000000000000;
mem[1864] = 80'h00000000000000000000;
mem[1865] = 80'h10100000010000010010;
mem[1866] = 80'h00109400000208004500;
mem[1867] = 80'h0010002e29940000fffd;
mem[1868] = 80'h00100fe6c0550102c000;
mem[1869] = 80'h00100001ffabffabffab;
mem[1870] = 80'h00106b1824b53418e8ec;
mem[1871] = 80'h0010992eb0c837a34d43;
mem[1872] = 80'h0110402a4425dcae21ef;
mem[1873] = 80'h00000000000000000000;
mem[1874] = 80'h00000000000000000000;
mem[1875] = 80'h00000000000000000000;
mem[1876] = 80'h10100000010000010010;
mem[1877] = 80'h00109400000208004500;
mem[1878] = 80'h0010002e29950000fffd;
mem[1879] = 80'h00100fe5c0550102c000;
mem[1880] = 80'h00100001ffabffabffab;
mem[1881] = 80'h00106a69fa99ec612a53;
mem[1882] = 80'h001052fc3725c2730412;
mem[1883] = 80'h011086b4aceb5f613a2c;
mem[1884] = 80'h00000000000000000000;
mem[1885] = 80'h00000000000000000000;
mem[1886] = 80'h00000000000000000000;
mem[1887] = 80'h10100000010000010010;
mem[1888] = 80'h00109400000208004500;
mem[1889] = 80'h0010002e29960000fffd;
mem[1890] = 80'h00100fe4c0550102c000;
mem[1891] = 80'h00100001ffabffabffab;
mem[1892] = 80'h001069fb98ec84eb6d93;
mem[1893] = 80'h00100e8bbf13dc034fe0;
mem[1894] = 80'h0110d5fd3b18189d0b52;
mem[1895] = 80'h00000000000000000000;
mem[1896] = 80'h10100000010000010010;
mem[1897] = 80'h00109400000208004500;
mem[1898] = 80'h0010002e29970000fffd;
mem[1899] = 80'h00100fe3c0550102c000;
mem[1900] = 80'h00100001ffabffabffab;
mem[1901] = 80'h0010688a46c05c92af2c;
mem[1902] = 80'h0010c55938fe29d310b1;
mem[1903] = 80'h0110bab6516321fc9ac5;
mem[1904] = 80'h00000000000000000000;
mem[1905] = 80'h00000000000000000000;
mem[1906] = 80'h00000000000000000000;
mem[1907] = 80'h00000000000000000000;
mem[1908] = 80'h10100000010000010010;
mem[1909] = 80'h00109400000208004500;
mem[1910] = 80'h0010002e29980000fffd;
mem[1911] = 80'h00100fe2c0550102c000;
mem[1912] = 80'h00100001ffabffabffab;
mem[1913] = 80'h001067b2113926c27292;
mem[1914] = 80'h00107f559dcba5c1a62b;
mem[1915] = 80'h0110d679ae37b23001bb;
mem[1916] = 80'h00000000000000000000;
mem[1917] = 80'h00000000000000000000;
mem[1918] = 80'h00000000000000000000;
mem[1919] = 80'h10100000010000010010;
mem[1920] = 80'h00109400000208004500;
mem[1921] = 80'h0010002e29990000fffd;
mem[1922] = 80'h00100fe1c0550102c000;
mem[1923] = 80'h00100001ffabffabffab;
mem[1924] = 80'h001066c3cf15febbb02d;
mem[1925] = 80'h0010b4871a265011e57a;
mem[1926] = 80'h0110ff2c17d6d4a516c2;
mem[1927] = 80'h00000000000000000000;
mem[1928] = 80'h10100000010000010010;
mem[1929] = 80'h00109400000208004500;
mem[1930] = 80'h0010002e299a0000fffd;
mem[1931] = 80'h00100fe0c0550102c000;
mem[1932] = 80'h00100001ffabffabffab;
mem[1933] = 80'h00106551ad609631f7ed;
mem[1934] = 80'h0010e8f092104e615788;
mem[1935] = 80'h0110053c3907e706d33d;
mem[1936] = 80'h00000000000000000000;
mem[1937] = 80'h00000000000000000000;
mem[1938] = 80'h00000000000000000000;
mem[1939] = 80'h10100000010000010010;
mem[1940] = 80'h00109400000208004500;
mem[1941] = 80'h0010002e299b0000fffd;
mem[1942] = 80'h00100fdfc0550102c000;
mem[1943] = 80'h00100001ffabffabffab;
mem[1944] = 80'h00106420734c4e483552;
mem[1945] = 80'h0010232215fdbbb0d9d9;
mem[1946] = 80'h01107b515afd6fcc0450;
mem[1947] = 80'h00000000000000000000;
mem[1948] = 80'h00000000000000000000;
mem[1949] = 80'h00000000000000000000;
mem[1950] = 80'h10100000010000010010;
mem[1951] = 80'h00109400000208004500;
mem[1952] = 80'h0010002e299c0000fffd;
mem[1953] = 80'h00100fdec0550102c000;
mem[1954] = 80'h00100001ffabffabffab;
mem[1955] = 80'h00106304b7a69f5cbad2;
mem[1956] = 80'h00109bcd04918751a33c;
mem[1957] = 80'h0110d99ce69bd0510b3a;
mem[1958] = 80'h00000000000000000000;
mem[1959] = 80'h00000000000000000000;
mem[1960] = 80'h00000000000000000000;
mem[1961] = 80'h10100000010000010010;
mem[1962] = 80'h00109400000208004500;
mem[1963] = 80'h0010002e299d0000fffd;
mem[1964] = 80'h00100fddc0550102c000;
mem[1965] = 80'h00100001ffabffabffab;
mem[1966] = 80'h00106275698a4725786d;
mem[1967] = 80'h0010501f837c7281b86d;
mem[1968] = 80'h011077dffe02ca6b2622;
mem[1969] = 80'h00000000000000000000;
mem[1970] = 80'h10100000010000010010;
mem[1971] = 80'h00109400000208004500;
mem[1972] = 80'h0010002e299e0000fffd;
mem[1973] = 80'h00100fdcc0550102c000;
mem[1974] = 80'h00100001ffabffabffab;
mem[1975] = 80'h001061e70bff2faf3fad;
mem[1976] = 80'h00100c680b4a6cf1339f;
mem[1977] = 80'h011032c237b8f88e0078;
mem[1978] = 80'h00000000000000000000;
mem[1979] = 80'h00000000000000000000;
mem[1980] = 80'h00000000000000000000;
mem[1981] = 80'h10100000010000010010;
mem[1982] = 80'h00109400000208004500;
mem[1983] = 80'h0010002e299f0000fffd;
mem[1984] = 80'h00100fdbc0550102c000;
mem[1985] = 80'h00100001ffabffabffab;
mem[1986] = 80'h00106096d5d3f7d6fd12;
mem[1987] = 80'h0010c7ba8ca79921bcce;
mem[1988] = 80'h011048aee1aa6e3c74db;
mem[1989] = 80'h00000000000000000000;
mem[1990] = 80'h00000000000000000000;
mem[1991] = 80'h00000000000000000000;
mem[1992] = 80'h10100000010000010010;
mem[1993] = 80'h00109400000208004500;
mem[1994] = 80'h0010002e29a00000fffd;
mem[1995] = 80'h00100fdac0550102c000;
mem[1996] = 80'h00100001ffabffabffab;
mem[1997] = 80'h00105fe5e843761fcc28;
mem[1998] = 80'h001073ff9047b71a6555;
mem[1999] = 80'h01101b8e39490fea85cb;
mem[2000] = 80'h00000000000000000000;
mem[2001] = 80'h00000000000000000000;
mem[2002] = 80'h00000000000000000000;
mem[2003] = 80'h10100000010000010010;
mem[2004] = 80'h00109400000208004500;
mem[2005] = 80'h0010002e29a10000fffd;
mem[2006] = 80'h00100fd9c0550102c000;
mem[2007] = 80'h00100001ffabffabffab;
mem[2008] = 80'h00105e94366fae660e97;
mem[2009] = 80'h0010b82d17aa42ca2604;
mem[2010] = 80'h011032db427dfeece7bd;
mem[2011] = 80'h00000000000000000000;
mem[2012] = 80'h10100000010000010010;
mem[2013] = 80'h00109400000208004500;
mem[2014] = 80'h0010002e29a20000fffd;
mem[2015] = 80'h00100fd8c0550102c000;
mem[2016] = 80'h00100001ffabffabffab;
mem[2017] = 80'h00105d06541ac6ec4957;
mem[2018] = 80'h0010e45a9f9c5cbae5f6;
mem[2019] = 80'h0110f3a3844e218e113b;
mem[2020] = 80'h00000000000000000000;
mem[2021] = 80'h00000000000000000000;
mem[2022] = 80'h00000000000000000000;
mem[2023] = 80'h00000000000000000000;
mem[2024] = 80'h10100000010000010010;
mem[2025] = 80'h00109400000208004500;
mem[2026] = 80'h0010002e29a30000fffd;
mem[2027] = 80'h00100fd7c0550102c000;
mem[2028] = 80'h00100001ffabffabffab;
mem[2029] = 80'h00105c778a361e958be8;
mem[2030] = 80'h00102f881871a96aa4a7;
mem[2031] = 80'h0110bc941c3455a04df3;
mem[2032] = 80'h00000000000000000000;
mem[2033] = 80'h00000000000000000000;
mem[2034] = 80'h00000000000000000000;
mem[2035] = 80'h10100000010000010010;
mem[2036] = 80'h00109400000208004500;
mem[2037] = 80'h0010002e29a40000fffd;
mem[2038] = 80'h00100fd6c0550102c000;
mem[2039] = 80'h00100001ffabffabffab;
mem[2040] = 80'h00105b534edccf810468;
mem[2041] = 80'h00109767091d958c0142;
mem[2042] = 80'h01109ed0abc22571cbaf;
mem[2043] = 80'h00000000000000000000;
mem[2044] = 80'h10100000010000010010;
mem[2045] = 80'h00109400000208004500;
mem[2046] = 80'h0010002e29a50000fffd;
mem[2047] = 80'h00100fd5c0550102c000;
mem[2048] = 80'h00100001ffabffabffab;
mem[2049] = 80'h00105a2290f017f8c6d7;
mem[2050] = 80'h00105cb58ef0605c4b13;
mem[2051] = 80'h01100d1d91eaa1430a82;
mem[2052] = 80'h00000000000000000000;
mem[2053] = 80'h00000000000000000000;
mem[2054] = 80'h00000000000000000000;
mem[2055] = 80'h10100000010000010010;
mem[2056] = 80'h00109400000208004500;
mem[2057] = 80'h0010002e29a60000fffd;
mem[2058] = 80'h00100fd4c0550102c000;
mem[2059] = 80'h00100001ffabffabffab;
mem[2060] = 80'h001059b0f2857f728117;
mem[2061] = 80'h001000c206c67e2c81e1;
mem[2062] = 80'h011076fd34acd78a83cc;
mem[2063] = 80'h00000000000000000000;
mem[2064] = 80'h00000000000000000000;
mem[2065] = 80'h00000000000000000000;
mem[2066] = 80'h10100000010000010010;
mem[2067] = 80'h00109400000208004500;
mem[2068] = 80'h0010002e29a70000fffd;
mem[2069] = 80'h00100fd3c0550102c000;
mem[2070] = 80'h00100001ffabffabffab;
mem[2071] = 80'h001058c12ca9a70b43a8;
mem[2072] = 80'h0010cb10812b8bfcffb0;
mem[2073] = 80'h01102c618b9607564525;
mem[2074] = 80'h00000000000000000000;
mem[2075] = 80'h00000000000000000000;
mem[2076] = 80'h00000000000000000000;
mem[2077] = 80'h10100000010000010010;
mem[2078] = 80'h00109400000208004500;
mem[2079] = 80'h0010002e29a80000fffd;
mem[2080] = 80'h00100fd2c0550102c000;
mem[2081] = 80'h00100001ffabffabffab;
mem[2082] = 80'h001057f97b50dd5b9e16;
mem[2083] = 80'h0010711c241e07ee0b2a;
mem[2084] = 80'h01102b00ddf0bb679d91;
mem[2085] = 80'h00000000000000000000;
mem[2086] = 80'h10100000010000010010;
mem[2087] = 80'h00109400000208004500;
mem[2088] = 80'h0010002e29a90000fffd;
mem[2089] = 80'h00100fd1c0550102c000;
mem[2090] = 80'h00100001ffabffabffab;
mem[2091] = 80'h00105688a57c05225ca9;
mem[2092] = 80'h0010bacea3f3f23e8a7b;
mem[2093] = 80'h01107263544fdc3ee6ac;
mem[2094] = 80'h00000000000000000000;
mem[2095] = 80'h00000000000000000000;
mem[2096] = 80'h00000000000000000000;
mem[2097] = 80'h10100000010000010010;
mem[2098] = 80'h00109400000208004500;
mem[2099] = 80'h0010002e29aa0000fffd;
mem[2100] = 80'h00100fd0c0550102c000;
mem[2101] = 80'h00100001ffabffabffab;
mem[2102] = 80'h0010551ac7096da81b69;
mem[2103] = 80'h0010e6b92bc5ec4e1f89;
mem[2104] = 80'h01101702257186e50cf4;
mem[2105] = 80'h00000000000000000000;
mem[2106] = 80'h00000000000000000000;
mem[2107] = 80'h00000000000000000000;
mem[2108] = 80'h10100000010000010010;
mem[2109] = 80'h00109400000208004500;
mem[2110] = 80'h0010002e29ab0000fffd;
mem[2111] = 80'h00100fcfc0550102c000;
mem[2112] = 80'h00100001ffabffabffab;
mem[2113] = 80'h0010546b1925b5d1d9d6;
mem[2114] = 80'h00102d6bac28199e16d8;
mem[2115] = 80'h0110dc501c6c4c564cd8;
mem[2116] = 80'h00000000000000000000;
mem[2117] = 80'h00000000000000000000;
mem[2118] = 80'h00000000000000000000;
mem[2119] = 80'h10100000010000010010;
mem[2120] = 80'h00109400000208004500;
mem[2121] = 80'h0010002e29ac0000fffd;
mem[2122] = 80'h00100fcec0550102c000;
mem[2123] = 80'h00100001ffabffabffab;
mem[2124] = 80'h0010534fddcf64c55656;
mem[2125] = 80'h00109584bd44257f6f3d;
mem[2126] = 80'h01102bce007179c22ecf;
mem[2127] = 80'h00000000000000000000;
mem[2128] = 80'h10100000010000010010;
mem[2129] = 80'h00109400000208004500;
mem[2130] = 80'h0010002e29ad0000fffd;
mem[2131] = 80'h00100fcdc0550102c000;
mem[2132] = 80'h00100001ffabffabffab;
mem[2133] = 80'h0010523e03e3bcbc94e9;
mem[2134] = 80'h00105e563aa9d0af176c;
mem[2135] = 80'h0110dbf4fb27d7d11957;
mem[2136] = 80'h00000000000000000000;
mem[2137] = 80'h00000000000000000000;
mem[2138] = 80'h00000000000000000000;
mem[2139] = 80'h00000000000000000000;
mem[2140] = 80'h10100000010000010010;
mem[2141] = 80'h00109400000208004500;
mem[2142] = 80'h0010002e29ae0000fffd;
mem[2143] = 80'h00100fccc0550102c000;
mem[2144] = 80'h00100001ffabffabffab;
mem[2145] = 80'h001051ac6196d436d329;
mem[2146] = 80'h00100221b29fcede5d9e;
mem[2147] = 80'h01108cbc3762c79aeeb1;
mem[2148] = 80'h00000000000000000000;
mem[2149] = 80'h00000000000000000000;
mem[2150] = 80'h00000000000000000000;
mem[2151] = 80'h10100000010000010010;
mem[2152] = 80'h00109400000208004500;
mem[2153] = 80'h0010002e29af0000fffd;
mem[2154] = 80'h00100fcbc0550102c000;
mem[2155] = 80'h00100001ffabffabffab;
mem[2156] = 80'h001050ddbfba0c4f1196;
mem[2157] = 80'h0010c9f335723b0e12cf;
mem[2158] = 80'h0110e084a3bae3be4ba4;
mem[2159] = 80'h00000000000000000000;
mem[2160] = 80'h10100000010000010010;
mem[2161] = 80'h00109400000208004500;
mem[2162] = 80'h0010002e29b00000fffd;
mem[2163] = 80'h00100fcac0550102c000;
mem[2164] = 80'h00100001ffabffabffab;
mem[2165] = 80'h00104fdcce6420976854;
mem[2166] = 80'h00107638f8f4d6fbbfaa;
mem[2167] = 80'h01105e84f47aec0193e6;
mem[2168] = 80'h00000000000000000000;
mem[2169] = 80'h00000000000000000000;
mem[2170] = 80'h00000000000000000000;
mem[2171] = 80'h10100000010000010010;
mem[2172] = 80'h00109400000208004500;
mem[2173] = 80'h0010002e29b10000fffd;
mem[2174] = 80'h00100fc9c0550102c000;
mem[2175] = 80'h00100001ffabffabffab;
mem[2176] = 80'h00104ead1048f8eeaaeb;
mem[2177] = 80'h0010bdea7f19232bfdfb;
mem[2178] = 80'h011044e05a244cb5b2cd;
mem[2179] = 80'h00000000000000000000;
mem[2180] = 80'h10100000010000010010;
mem[2181] = 80'h00109400000208004500;
mem[2182] = 80'h0010002e29b20000fffd;
mem[2183] = 80'h00100fc8c0550102c000;
mem[2184] = 80'h00100001ffabffabffab;
mem[2185] = 80'h00104d3f723d9064ed2b;
mem[2186] = 80'h0010e19df72f3d5bbf09;
mem[2187] = 80'h0110ad31408e2350d989;
mem[2188] = 80'h00000000000000000000;
mem[2189] = 80'h00000000000000000000;
mem[2190] = 80'h00000000000000000000;
mem[2191] = 80'h00000000000000000000;
mem[2192] = 80'h10100000010000010010;
mem[2193] = 80'h00109400000208004500;
mem[2194] = 80'h0010002e29b30000fffd;
mem[2195] = 80'h00100fc7c0550102c000;
mem[2196] = 80'h00100001ffabffabffab;
mem[2197] = 80'h00104c4eac11481d2f94;
mem[2198] = 80'h00102a4f70c2c88bc058;
mem[2199] = 80'h0110c49ca75b0e0ee6e4;
mem[2200] = 80'h00000000000000000000;
mem[2201] = 80'h00000000000000000000;
mem[2202] = 80'h00000000000000000000;
mem[2203] = 80'h10100000010000010010;
mem[2204] = 80'h00109400000208004500;
mem[2205] = 80'h0010002e29b40000fffd;
mem[2206] = 80'h00100fc6c0550102c000;
mem[2207] = 80'h00100001ffabffabffab;
mem[2208] = 80'h00104b6a68fb9909a014;
mem[2209] = 80'h001092a061aef46abbbd;
mem[2210] = 80'h0110556018a4dfe07c20;
mem[2211] = 80'h00000000000000000000;
mem[2212] = 80'h00000000000000000000;
mem[2213] = 80'h00000000000000000000;
mem[2214] = 80'h10100000010000010010;
mem[2215] = 80'h00109400000208004500;
mem[2216] = 80'h0010002e29b50000fffd;
mem[2217] = 80'h00100fc5c0550102c000;
mem[2218] = 80'h00100001ffabffabffab;
mem[2219] = 80'h00104a1bb6d7417062ab;
mem[2220] = 80'h00105972e64301bab0ec;
mem[2221] = 80'h0110f8507043748407e7;
mem[2222] = 80'h00000000000000000000;
mem[2223] = 80'h10100000010000010010;
mem[2224] = 80'h00109400000208004500;
mem[2225] = 80'h0010002e29b60000fffd;
mem[2226] = 80'h00100fc4c0550102c000;
mem[2227] = 80'h00100001ffabffabffab;
mem[2228] = 80'h00104989d4a229fa256b;
mem[2229] = 80'h001005056e751fca3b1e;
mem[2230] = 80'h0110bd4d06be0207c436;
mem[2231] = 80'h00000000000000000000;
mem[2232] = 80'h00000000000000000000;
mem[2233] = 80'h00000000000000000000;
mem[2234] = 80'h10100000010000010010;
mem[2235] = 80'h00109400000208004500;
mem[2236] = 80'h0010002e29b70000fffd;
mem[2237] = 80'h00100fc3c0550102c000;
mem[2238] = 80'h00100001ffabffabffab;
mem[2239] = 80'h001048f80a8ef183e7d4;
mem[2240] = 80'h0010ced7e998ea19a44f;
mem[2241] = 80'h01109d02ef43386f5e51;
mem[2242] = 80'h00000000000000000000;
mem[2243] = 80'h00000000000000000000;
mem[2244] = 80'h00000000000000000000;
mem[2245] = 80'h10100000010000010010;
mem[2246] = 80'h00109400000208004500;
mem[2247] = 80'h0010002e29b80000fffd;
mem[2248] = 80'h00100fc2c0550102c000;
mem[2249] = 80'h00100001ffabffabffab;
mem[2250] = 80'h001047c05d778bd33a6a;
mem[2251] = 80'h001074db4cad660b51d5;
mem[2252] = 80'h0110a95271ce7f3316dd;
mem[2253] = 80'h00000000000000000000;
mem[2254] = 80'h00000000000000000000;
mem[2255] = 80'h00000000000000000000;
mem[2256] = 80'h10100000010000010010;
mem[2257] = 80'h00109400000208004500;
mem[2258] = 80'h0010002e29b90000fffd;
mem[2259] = 80'h00100fc1c0550102c000;
mem[2260] = 80'h00100001ffabffabffab;
mem[2261] = 80'h001046b1835b53aaf8d5;
mem[2262] = 80'h0010bf09cb4093db5184;
mem[2263] = 80'h0110d898a12fb5d60461;
mem[2264] = 80'h00000000000000000000;
mem[2265] = 80'h00000000000000000000;
mem[2266] = 80'h00000000000000000000;
mem[2267] = 80'h10100000010000010010;
mem[2268] = 80'h00109400000208004500;
mem[2269] = 80'h0010002e29ba0000fffd;
mem[2270] = 80'h00100fc0c0550102c000;
mem[2271] = 80'h00100001ffabffabffab;
mem[2272] = 80'h00104523e12e3b20bf15;
mem[2273] = 80'h0010e37e43768dabe276;
mem[2274] = 80'h011011b936a76a821ab5;
mem[2275] = 80'h00000000000000000000;
mem[2276] = 80'h10100000010000010010;
mem[2277] = 80'h00109400000208004500;
mem[2278] = 80'h0010002e29bb0000fffd;
mem[2279] = 80'h00100fbfc0550102c000;
mem[2280] = 80'h00100001ffabffabffab;
mem[2281] = 80'h001044523f02e3597daa;
mem[2282] = 80'h001028acc49b787bac27;
mem[2283] = 80'h01104eb0bb0b8bcb6f9e;
mem[2284] = 80'h00000000000000000000;
mem[2285] = 80'h00000000000000000000;
mem[2286] = 80'h00000000000000000000;
mem[2287] = 80'h10100000010000010010;
mem[2288] = 80'h00109400000208004500;
mem[2289] = 80'h0010002e29bc0000fffd;
mem[2290] = 80'h00100fbec0550102c000;
mem[2291] = 80'h00100001ffabffabffab;
mem[2292] = 80'h00104376fbe8324df22a;
mem[2293] = 80'h00109043d5f7449a16c2;
mem[2294] = 80'h0110fa29e0660c7aa27d;
mem[2295] = 80'h00000000000000000000;
mem[2296] = 80'h00000000000000000000;
mem[2297] = 80'h00000000000000000000;
mem[2298] = 80'h10100000010000010010;
mem[2299] = 80'h00109400000208004500;
mem[2300] = 80'h0010002e29bd0000fffd;
mem[2301] = 80'h00100fbdc0550102c000;
mem[2302] = 80'h00100001ffabffabffab;
mem[2303] = 80'h0010420725c4ea343095;
mem[2304] = 80'h00105b91521ab14a4c93;
mem[2305] = 80'h01106a976749a276b8d8;
mem[2306] = 80'h00000000000000000000;
mem[2307] = 80'h00000000000000000000;
mem[2308] = 80'h00000000000000000000;
mem[2309] = 80'h10100000010000010010;
mem[2310] = 80'h00109400000208004500;
mem[2311] = 80'h0010002e29be0000fffd;
mem[2312] = 80'h00100fbcc0550102c000;
mem[2313] = 80'h00100001ffabffabffab;
mem[2314] = 80'h0010419547b182be7755;
mem[2315] = 80'h001007e6da2caf3a8961;
mem[2316] = 80'h0110014960adab8e62bd;
mem[2317] = 80'h00000000000000000000;
mem[2318] = 80'h10100000010000010010;
mem[2319] = 80'h00109400000208004500;
mem[2320] = 80'h0010002e29bf0000fffd;
mem[2321] = 80'h00100fbbc0550102c000;
mem[2322] = 80'h00100001ffabffabffab;
mem[2323] = 80'h001040e4999d5ac7b5ea;
mem[2324] = 80'h0010cc345dc15aeac830;
mem[2325] = 80'h01104e7e793c20933baa;
mem[2326] = 80'h00000000000000000000;
mem[2327] = 80'h00000000000000000000;
mem[2328] = 80'h00000000000000000000;
mem[2329] = 80'h10100000010000010010;
mem[2330] = 80'h00109400000208004500;
mem[2331] = 80'h0010002e29c00000fffd;
mem[2332] = 80'h00100fbac0550102c000;
mem[2333] = 80'h00100001ffabffabffab;
mem[2334] = 80'h00103f733c90812c1520;
mem[2335] = 80'h00106f6ce3ecf34d3857;
mem[2336] = 80'h0110c16bad45afe10aa6;
mem[2337] = 80'h00000000000000000000;
mem[2338] = 80'h00000000000000000000;
mem[2339] = 80'h00000000000000000000;
mem[2340] = 80'h10100000010000010010;
mem[2341] = 80'h00109400000208004500;
mem[2342] = 80'h0010002e29c10000fffd;
mem[2343] = 80'h00100fb9c0550102c000;
mem[2344] = 80'h00100001ffabffabffab;
mem[2345] = 80'h00103e02e2bc5955d79f;
mem[2346] = 80'h0010a4be6401069cb906;
mem[2347] = 80'h0110af3836b0a94e6c9a;
mem[2348] = 80'h00000000000000000000;
mem[2349] = 80'h00000000000000000000;
mem[2350] = 80'h00000000000000000000;
mem[2351] = 80'h10100000010000010010;
mem[2352] = 80'h00109400000208004500;
mem[2353] = 80'h0010002e29c20000fffd;
mem[2354] = 80'h00100fb8c0550102c000;
mem[2355] = 80'h00100001ffabffabffab;
mem[2356] = 80'h00103d9080c931df905f;
mem[2357] = 80'h0010f8c9ec3718ec3cf4;
mem[2358] = 80'h0110c92a7b5abd811f77;
mem[2359] = 80'h00000000000000000000;
mem[2360] = 80'h10100000010000010010;
mem[2361] = 80'h00109400000208004500;
mem[2362] = 80'h0010002e29c30000fffd;
mem[2363] = 80'h00100fb7c0550102c000;
mem[2364] = 80'h00100001ffabffabffab;
mem[2365] = 80'h00103ce15ee5e9a652e0;
mem[2366] = 80'h0010331b6bdaed3c24a5;
mem[2367] = 80'h0110323a44a050d62e37;
mem[2368] = 80'h00000000000000000000;
mem[2369] = 80'h00000000000000000000;
mem[2370] = 80'h00000000000000000000;
mem[2371] = 80'h10100000010000010010;
mem[2372] = 80'h00109400000208004500;
mem[2373] = 80'h0010002e29c40000fffd;
mem[2374] = 80'h00100fb6c0550102c000;
mem[2375] = 80'h00100001ffabffabffab;
mem[2376] = 80'h00103bc59a0f38b2dd60;
mem[2377] = 80'h00108bf47ab6d1dd5c40;
mem[2378] = 80'h0110f695e8b81f1388b8;
mem[2379] = 80'h00000000000000000000;
mem[2380] = 80'h00000000000000000000;
mem[2381] = 80'h00000000000000000000;
mem[2382] = 80'h10100000010000010010;
mem[2383] = 80'h00109400000208004500;
mem[2384] = 80'h0010002e29c50000fffd;
mem[2385] = 80'h00100fb5c0550102c000;
mem[2386] = 80'h00100001ffabffabffab;
mem[2387] = 80'h00103ab44423e0cb1fdf;
mem[2388] = 80'h00104026fd5b240dd511;
mem[2389] = 80'h0110265f237deee2c75d;
mem[2390] = 80'h00000000000000000000;
mem[2391] = 80'h10100000010000010010;
mem[2392] = 80'h00109400000208004500;
mem[2393] = 80'h0010002e29c60000fffd;
mem[2394] = 80'h00100fb4c0550102c000;
mem[2395] = 80'h00100001ffabffabffab;
mem[2396] = 80'h0010392626568841581f;
mem[2397] = 80'h00101c51756d3a7d5fe3;
mem[2398] = 80'h01105073439066cf4081;
mem[2399] = 80'h00000000000000000000;
mem[2400] = 80'h00000000000000000000;
mem[2401] = 80'h00000000000000000000;
mem[2402] = 80'h00000000000000000000;
mem[2403] = 80'h10100000010000010010;
mem[2404] = 80'h00109400000208004500;
mem[2405] = 80'h0010002e29c70000fffd;
mem[2406] = 80'h00100fb3c0550102c000;
mem[2407] = 80'h00100001ffabffabffab;
mem[2408] = 80'h00103857f87a50389aa0;
mem[2409] = 80'h0010d783f280cfad21b2;
mem[2410] = 80'h01100aef1e01b8f8ca45;
mem[2411] = 80'h00000000000000000000;
mem[2412] = 80'h00000000000000000000;
mem[2413] = 80'h00000000000000000000;
mem[2414] = 80'h10100000010000010010;
mem[2415] = 80'h00109400000208004500;
mem[2416] = 80'h0010002e29c80000fffd;
mem[2417] = 80'h00100fb2c0550102c000;
mem[2418] = 80'h00100001ffabffabffab;
mem[2419] = 80'h0010376faf832a68471e;
mem[2420] = 80'h00106d8f57b543bf9628;
mem[2421] = 80'h01105511b348696cb1dc;
mem[2422] = 80'h00000000000000000000;
mem[2423] = 80'h10100000010000010010;
mem[2424] = 80'h00109400000208004500;
mem[2425] = 80'h0010002e29c90000fffd;
mem[2426] = 80'h00100fb1c0550102c000;
mem[2427] = 80'h00100001ffabffabffab;
mem[2428] = 80'h0010361e71aff21185a1;
mem[2429] = 80'h0010a65dd058b66fd579;
mem[2430] = 80'h01107c44619a752a7f9c;
mem[2431] = 80'h00000000000000000000;
mem[2432] = 80'h00000000000000000000;
mem[2433] = 80'h00000000000000000000;
mem[2434] = 80'h10100000010000010010;
mem[2435] = 80'h00109400000208004500;
mem[2436] = 80'h0010002e29ca0000fffd;
mem[2437] = 80'h00100fb0c0550102c000;
mem[2438] = 80'h00100001ffabffabffab;
mem[2439] = 80'h0010358c13da9a9bc261;
mem[2440] = 80'h0010fa2a586ea810868b;
mem[2441] = 80'h011089e64e80d921fec3;
mem[2442] = 80'h00000000000000000000;
mem[2443] = 80'h00000000000000000000;
mem[2444] = 80'h00000000000000000000;
mem[2445] = 80'h10100000010000010010;
mem[2446] = 80'h00109400000208004500;
mem[2447] = 80'h0010002e29cb0000fffd;
mem[2448] = 80'h00100fafc0550102c000;
mem[2449] = 80'h00100001ffabffabffab;
mem[2450] = 80'h001034fdcdf642e200de;
mem[2451] = 80'h001031f8df835dc0c9da;
mem[2452] = 80'h0110e5de9a550bd32cdd;
mem[2453] = 80'h00000000000000000000;
mem[2454] = 80'h10100000010000010010;
mem[2455] = 80'h00109400000208004500;
mem[2456] = 80'h0010002e29cc0000fffd;
mem[2457] = 80'h00100faec0550102c000;
mem[2458] = 80'h00100001ffabffabffab;
mem[2459] = 80'h001033d9091c93f68f5e;
mem[2460] = 80'h00108917ceef6121f23f;
mem[2461] = 80'h011079ee7a5ed1f7c2fb;
mem[2462] = 80'h00000000000000000000;
mem[2463] = 80'h00000000000000000000;
mem[2464] = 80'h00000000000000000000;
mem[2465] = 80'h00000000000000000000;
mem[2466] = 80'h10100000010000010010;
mem[2467] = 80'h00109400000208004500;
mem[2468] = 80'h0010002e29cd0000fffd;
mem[2469] = 80'h00100fadc0550102c000;
mem[2470] = 80'h00100001ffabffabffab;
mem[2471] = 80'h001032a8d7304b8f4de1;
mem[2472] = 80'h001042c5490294f1896e;
mem[2473] = 80'h0110dc87d6063c1f0a65;
mem[2474] = 80'h00000000000000000000;
mem[2475] = 80'h00000000000000000000;
mem[2476] = 80'h00000000000000000000;
mem[2477] = 80'h10100000010000010010;
mem[2478] = 80'h00109400000208004500;
mem[2479] = 80'h0010002e29ce0000fffd;
mem[2480] = 80'h00100facc0550102c000;
mem[2481] = 80'h00100001ffabffabffab;
mem[2482] = 80'h0010313ab54523050a21;
mem[2483] = 80'h00101eb2c1348a810d9c;
mem[2484] = 80'h011089a4eab00d8eebd0;
mem[2485] = 80'h00000000000000000000;
mem[2486] = 80'h10100000010000010010;
mem[2487] = 80'h00109400000208004500;
mem[2488] = 80'h0010002e29cf0000fffd;
mem[2489] = 80'h00100fabc0550102c000;
mem[2490] = 80'h00100001ffabffabffab;
mem[2491] = 80'h0010304b6b69fb7cc89e;
mem[2492] = 80'h0010d56046d97f518dcd;
mem[2493] = 80'h0110e3f692dfad8d15e2;
mem[2494] = 80'h00000000000000000000;
mem[2495] = 80'h00000000000000000000;
mem[2496] = 80'h00000000000000000000;
mem[2497] = 80'h10100000010000010010;
mem[2498] = 80'h00109400000208004500;
mem[2499] = 80'h0010002e29d00000fffd;
mem[2500] = 80'h00100faac0550102c000;
mem[2501] = 80'h00100001ffabffabffab;
mem[2502] = 80'h00102f4a1ab7d7a4b15c;
mem[2503] = 80'h00106aab8b5f92a462a8;
mem[2504] = 80'h011036580b4db553800d;
mem[2505] = 80'h00000000000000000000;
mem[2506] = 80'h00000000000000000000;
mem[2507] = 80'h00000000000000000000;
mem[2508] = 80'h00000000000000000000;
mem[2509] = 80'h10100000010000010010;
mem[2510] = 80'h00109400000208004500;
mem[2511] = 80'h0010002e29d10000fffd;
mem[2512] = 80'h00100fa9c0550102c000;
mem[2513] = 80'h00100001ffabffabffab;
mem[2514] = 80'h00102e3bc49b0fdd73e3;
mem[2515] = 80'h0010a1790cb2677463f9;
mem[2516] = 80'h011074a39b2bb4e45c3e;
mem[2517] = 80'h00000000000000000000;
mem[2518] = 80'h10100000010000010010;
mem[2519] = 80'h00109400000208004500;
mem[2520] = 80'h0010002e29d20000fffd;
mem[2521] = 80'h00100fa8c0550102c000;
mem[2522] = 80'h00100001ffabffabffab;
mem[2523] = 80'h00102da9a6ee67573423;
mem[2524] = 80'h0010fd0e84847904e10b;
mem[2525] = 80'h01108b26292365651e2b;
mem[2526] = 80'h00000000000000000000;
mem[2527] = 80'h00000000000000000000;
mem[2528] = 80'h00000000000000000000;
mem[2529] = 80'h10100000010000010010;
mem[2530] = 80'h00109400000208004500;
mem[2531] = 80'h0010002e29d30000fffd;
mem[2532] = 80'h00100fa7c0550102c000;
mem[2533] = 80'h00100001ffabffabffab;
mem[2534] = 80'h00102cd878c2bf2ef69c;
mem[2535] = 80'h001036dc03698cd49f5a;
mem[2536] = 80'h0110d1ba6c6a0131c22f;
mem[2537] = 80'h00000000000000000000;
mem[2538] = 80'h00000000000000000000;
mem[2539] = 80'h00000000000000000000;
mem[2540] = 80'h10100000010000010010;
mem[2541] = 80'h00109400000208004500;
mem[2542] = 80'h0010002e29d40000fffd;
mem[2543] = 80'h00100fa6c0550102c000;
mem[2544] = 80'h00100001ffabffabffab;
mem[2545] = 80'h00102bfcbc286e3a791c;
mem[2546] = 80'h00108e331205b03426bf;
mem[2547] = 80'h01100740b21707cf116c;
mem[2548] = 80'h00000000000000000000;
mem[2549] = 80'h10100000010000010010;
mem[2550] = 80'h00109400000208004500;
mem[2551] = 80'h0010002e29d50000fffd;
mem[2552] = 80'h00100fa5c0550102c000;
mem[2553] = 80'h00100001ffabffabffab;
mem[2554] = 80'h00102a8d6204b643bba3;
mem[2555] = 80'h001045e195e845e46fee;
mem[2556] = 80'h0110c1deae0bc59707b7;
mem[2557] = 80'h00000000000000000000;
mem[2558] = 80'h00000000000000000000;
mem[2559] = 80'h00000000000000000000;
mem[2560] = 80'h00000000000000000000;
mem[2561] = 80'h10100000010000010010;
mem[2562] = 80'h00109400000208004500;
mem[2563] = 80'h0010002e29d60000fffd;
mem[2564] = 80'h00100fa4c0550102c000;
mem[2565] = 80'h00100001ffabffabffab;
mem[2566] = 80'h0010291f0071dec9fc63;
mem[2567] = 80'h001019961dde5b94ba1c;
mem[2568] = 80'h0110a97304a9b1321f11;
mem[2569] = 80'h00000000000000000000;
mem[2570] = 80'h00000000000000000000;
mem[2571] = 80'h00000000000000000000;
mem[2572] = 80'h10100000010000010010;
mem[2573] = 80'h00109400000208004500;
mem[2574] = 80'h0010002e29d70000fffd;
mem[2575] = 80'h00100fa3c0550102c000;
mem[2576] = 80'h00100001ffabffabffab;
mem[2577] = 80'h0010286ede5d06b03edc;
mem[2578] = 80'h0010d2449a33ae44fb4d;
mem[2579] = 80'h0110e644b7579007a38f;
mem[2580] = 80'h00000000000000000000;
mem[2581] = 80'h10100000010000010010;
mem[2582] = 80'h00109400000208004500;
mem[2583] = 80'h0010002e29d80000fffd;
mem[2584] = 80'h00100fa2c0550102c000;
mem[2585] = 80'h00100001ffabffabffab;
mem[2586] = 80'h0010275689a47ce0e362;
mem[2587] = 80'h001068483f062256cfd7;
mem[2588] = 80'h0110f7715dd357c42032;
mem[2589] = 80'h00000000000000000000;
mem[2590] = 80'h00000000000000000000;
mem[2591] = 80'h00000000000000000000;
mem[2592] = 80'h00000000000000000000;
mem[2593] = 80'h10100000010000010010;
mem[2594] = 80'h00109400000208004500;
mem[2595] = 80'h0010002e29d90000fffd;
mem[2596] = 80'h00100fa1c0550102c000;
mem[2597] = 80'h00100001ffabffabffab;
mem[2598] = 80'h001026275788a49921dd;
mem[2599] = 80'h0010a39ab8ebd7868f86;
mem[2600] = 80'h01108b776cce92e0db18;
mem[2601] = 80'h00000000000000000000;
mem[2602] = 80'h10100000010000010010;
mem[2603] = 80'h00109400000208004500;
mem[2604] = 80'h0010002e29da0000fffd;
mem[2605] = 80'h00100fa0c0550102c000;
mem[2606] = 80'h00100001ffabffabffab;
mem[2607] = 80'h001025b535fdcc13661d;
mem[2608] = 80'h0010ffed30ddc9f63b74;
mem[2609] = 80'h0110dbc160240bd7ddd8;
mem[2610] = 80'h00000000000000000000;
mem[2611] = 80'h00000000000000000000;
mem[2612] = 80'h00000000000000000000;
mem[2613] = 80'h00000000000000000000;
mem[2614] = 80'h10100000010000010010;
mem[2615] = 80'h00109400000208004500;
mem[2616] = 80'h0010002e29db0000fffd;
mem[2617] = 80'h00100f9fc0550102c000;
mem[2618] = 80'h00100001ffabffabffab;
mem[2619] = 80'h001024c4ebd1146aa4a2;
mem[2620] = 80'h0010343fb7303c263325;
mem[2621] = 80'h011023a2b7fffd5ef8d5;
mem[2622] = 80'h00000000000000000000;
mem[2623] = 80'h00000000000000000000;
mem[2624] = 80'h00000000000000000000;
mem[2625] = 80'h10100000010000010010;
mem[2626] = 80'h00109400000208004500;
mem[2627] = 80'h0010002e29dc0000fffd;
mem[2628] = 80'h00100f9ec0550102c000;
mem[2629] = 80'h00100001ffabffabffab;
mem[2630] = 80'h001023e02f3bc57e2b22;
mem[2631] = 80'h00108cd0a65c00c74ac0;
mem[2632] = 80'h0110d43c695288cc37f0;
mem[2633] = 80'h00000000000000000000;
mem[2634] = 80'h10100000010000010010;
mem[2635] = 80'h00109400000208004500;
mem[2636] = 80'h0010002e29dd0000fffd;
mem[2637] = 80'h00100f9dc0550102c000;
mem[2638] = 80'h00100001ffabffabffab;
mem[2639] = 80'h00102291f1171d07e99d;
mem[2640] = 80'h0010470221b1f514d391;
mem[2641] = 80'h01105ed5558291a1dd8f;
mem[2642] = 80'h00000000000000000000;
mem[2643] = 80'h00000000000000000000;
mem[2644] = 80'h00000000000000000000;
mem[2645] = 80'h00000000000000000000;
mem[2646] = 80'h10100000010000010010;
mem[2647] = 80'h00109400000208004500;
mem[2648] = 80'h0010002e29de0000fffd;
mem[2649] = 80'h00100f9cc0550102c000;
mem[2650] = 80'h00100001ffabffabffab;
mem[2651] = 80'h001021039362758dae5d;
mem[2652] = 80'h00101b75a987eb645863;
mem[2653] = 80'h01101bc803220c2b40de;
mem[2654] = 80'h00000000000000000000;
mem[2655] = 80'h00000000000000000000;
mem[2656] = 80'h00000000000000000000;
mem[2657] = 80'h10100000010000010010;
mem[2658] = 80'h00109400000208004500;
mem[2659] = 80'h0010002e29df0000fffd;
mem[2660] = 80'h00100f9bc0550102c000;
mem[2661] = 80'h00100001ffabffabffab;
mem[2662] = 80'h001020724d4eadf46ce2;
mem[2663] = 80'h0010d0a72e6a1eb45732;
mem[2664] = 80'h01107a3c883337c68081;
mem[2665] = 80'h00000000000000000000;
mem[2666] = 80'h10100000010000010010;
mem[2667] = 80'h00109400000208004500;
mem[2668] = 80'h0010002e29e00000fffd;
mem[2669] = 80'h00100f9ac0550102c000;
mem[2670] = 80'h00100001ffabffabffab;
mem[2671] = 80'h00101f0170de2c3d5dd8;
mem[2672] = 80'h001064e2328a308f8ea9;
mem[2673] = 80'h0110291c6649c3aabe91;
mem[2674] = 80'h00000000000000000000;
mem[2675] = 80'h00000000000000000000;
mem[2676] = 80'h00000000000000000000;
mem[2677] = 80'h10100000010000010010;
mem[2678] = 80'h00109400000208004500;
mem[2679] = 80'h0010002e29e10000fffd;
mem[2680] = 80'h00100f99c0550102c000;
mem[2681] = 80'h00100001ffabffabffab;
mem[2682] = 80'h00101e70aef2f4449f67;
mem[2683] = 80'h0010af30b567c55fcdf8;
mem[2684] = 80'h01100049a6b679c05bec;
mem[2685] = 80'h00000000000000000000;
mem[2686] = 80'h00000000000000000000;
mem[2687] = 80'h00000000000000000000;
mem[2688] = 80'h10100000010000010010;
mem[2689] = 80'h00109400000208004500;
mem[2690] = 80'h0010002e29e20000fffd;
mem[2691] = 80'h00100f98c0550102c000;
mem[2692] = 80'h00100001ffabffabffab;
mem[2693] = 80'h00101de2cc879cced8a7;
mem[2694] = 80'h0010f3473d51db2f8e0a;
mem[2695] = 80'h0110daa92ba20dac82b6;
mem[2696] = 80'h00000000000000000000;
mem[2697] = 80'h00000000000000000000;
mem[2698] = 80'h00000000000000000000;
mem[2699] = 80'h10100000010000010010;
mem[2700] = 80'h00109400000208004500;
mem[2701] = 80'h0010002e29e30000fffd;
mem[2702] = 80'h00100f97c0550102c000;
mem[2703] = 80'h00100001ffabffabffab;
mem[2704] = 80'h00101c9312ab44b71a18;
mem[2705] = 80'h00103895babc2effd15b;
mem[2706] = 80'h0110b5e2c8623725a45d;
mem[2707] = 80'h00000000000000000000;
mem[2708] = 80'h10100000010000010010;
mem[2709] = 80'h00109400000208004500;
mem[2710] = 80'h0010002e29e40000fffd;
mem[2711] = 80'h00100f96c0550102c000;
mem[2712] = 80'h00100001ffabffabffab;
mem[2713] = 80'h00101bb7d64195a39598;
mem[2714] = 80'h0010807aabd0121ee9be;
mem[2715] = 80'h01107c813e214f60680b;
mem[2716] = 80'h00000000000000000000;
mem[2717] = 80'h00000000000000000000;
mem[2718] = 80'h00000000000000000000;
mem[2719] = 80'h10100000010000010010;
mem[2720] = 80'h00109400000208004500;
mem[2721] = 80'h0010002e29e50000fffd;
mem[2722] = 80'h00100f95c0550102c000;
mem[2723] = 80'h00100001ffabffabffab;
mem[2724] = 80'h00101ac6086d4dda5727;
mem[2725] = 80'h00104ba82c3de7cea1ef;
mem[2726] = 80'h0110892eacf83ab01b92;
mem[2727] = 80'h00000000000000000000;
mem[2728] = 80'h00000000000000000000;
mem[2729] = 80'h00000000000000000000;
mem[2730] = 80'h10100000010000010010;
mem[2731] = 80'h00109400000208004500;
mem[2732] = 80'h0010002e29e60000fffd;
mem[2733] = 80'h00100f94c0550102c000;
mem[2734] = 80'h00100001ffabffabffab;
mem[2735] = 80'h001019546a18255010e7;
mem[2736] = 80'h001017dfa40bf9be151d;
mem[2737] = 80'h0110d998a1fc9d79b40c;
mem[2738] = 80'h00000000000000000000;
mem[2739] = 80'h00000000000000000000;
mem[2740] = 80'h00000000000000000000;
mem[2741] = 80'h10100000010000010010;
mem[2742] = 80'h00109400000208004500;
mem[2743] = 80'h0010002e29e70000fffd;
mem[2744] = 80'h00100f93c0550102c000;
mem[2745] = 80'h00100001ffabffabffab;
mem[2746] = 80'h00101825b434fd29d258;
mem[2747] = 80'h0010dc0d23e60c6f964c;
mem[2748] = 80'h0110d1a9efc94960b5c7;
mem[2749] = 80'h00000000000000000000;
mem[2750] = 80'h10100000010000010010;
mem[2751] = 80'h00109400000208004500;
mem[2752] = 80'h0010002e29e80000fffd;
mem[2753] = 80'h00100f92c0550102c000;
mem[2754] = 80'h00100001ffabffabffab;
mem[2755] = 80'h0010171de3cd87790fe6;
mem[2756] = 80'h0010660186d3807d60d6;
mem[2757] = 80'h0110b0aaeee16be0250f;
mem[2758] = 80'h00000000000000000000;
mem[2759] = 80'h00000000000000000000;
mem[2760] = 80'h00000000000000000000;
mem[2761] = 80'h00000000000000000000;
mem[2762] = 80'h10100000010000010010;
mem[2763] = 80'h00109400000208004500;
mem[2764] = 80'h0010002e29e90000fffd;
mem[2765] = 80'h00100f91c0550102c000;
mem[2766] = 80'h00100001ffabffabffab;
mem[2767] = 80'h0010166c3de15f00cd59;
mem[2768] = 80'h0010add3013e75ad6187;
mem[2769] = 80'h0110f25106c0a770a733;
mem[2770] = 80'h00000000000000000000;
mem[2771] = 80'h00000000000000000000;
mem[2772] = 80'h00000000000000000000;
mem[2773] = 80'h10100000010000010010;
mem[2774] = 80'h00109400000208004500;
mem[2775] = 80'h0010002e29ea0000fffd;
mem[2776] = 80'h00100f90c0550102c000;
mem[2777] = 80'h00100001ffabffabffab;
mem[2778] = 80'h001015fe5f94378a8a99;
mem[2779] = 80'h0010f1a489086bddf475;
mem[2780] = 80'h01109730561853f9bbae;
mem[2781] = 80'h00000000000000000000;
mem[2782] = 80'h10100000010000010010;
mem[2783] = 80'h00109400000208004500;
mem[2784] = 80'h0010002e29eb0000fffd;
mem[2785] = 80'h00100f8fc0550102c000;
mem[2786] = 80'h00100001ffabffabffab;
mem[2787] = 80'h0010148f81b8eff34826;
mem[2788] = 80'h00103a760ee59e0d7d24;
mem[2789] = 80'h011047fa85162f3d7cc8;
mem[2790] = 80'h00000000000000000000;
mem[2791] = 80'h00000000000000000000;
mem[2792] = 80'h00000000000000000000;
mem[2793] = 80'h10100000010000010010;
mem[2794] = 80'h00109400000208004500;
mem[2795] = 80'h0010002e29ec0000fffd;
mem[2796] = 80'h00100f8ec0550102c000;
mem[2797] = 80'h00100001ffabffabffab;
mem[2798] = 80'h001013ab45523ee7c7a6;
mem[2799] = 80'h001082991f89a2ec04c1;
mem[2800] = 80'h0110b064a63f937774a6;
mem[2801] = 80'h00000000000000000000;
mem[2802] = 80'h10100000010000010010;
mem[2803] = 80'h00109400000208004500;
mem[2804] = 80'h0010002e29ed0000fffd;
mem[2805] = 80'h00100f8dc0550102c000;
mem[2806] = 80'h00100001ffabffabffab;
mem[2807] = 80'h001012da9b7ee69e0519;
mem[2808] = 80'h0010494b9864573c7c90;
mem[2809] = 80'h0110405e70145333dd30;
mem[2810] = 80'h00000000000000000000;
mem[2811] = 80'h00000000000000000000;
mem[2812] = 80'h00000000000000000000;
mem[2813] = 80'h00000000000000000000;
mem[2814] = 80'h10100000010000010010;
mem[2815] = 80'h00109400000208004500;
mem[2816] = 80'h0010002e29ee0000fffd;
mem[2817] = 80'h00100f8cc0550102c000;
mem[2818] = 80'h00100001ffabffabffab;
mem[2819] = 80'h00101148f90b8e1442d9;
mem[2820] = 80'h0010153c1052494cb862;
mem[2821] = 80'h011018b1e4cff33466b5;
mem[2822] = 80'h00000000000000000000;
mem[2823] = 80'h00000000000000000000;
mem[2824] = 80'h00000000000000000000;
mem[2825] = 80'h10100000010000010010;
mem[2826] = 80'h00109400000208004500;
mem[2827] = 80'h0010002e29ef0000fffd;
mem[2828] = 80'h00100f8bc0550102c000;
mem[2829] = 80'h00100001ffabffabffab;
mem[2830] = 80'h001010392727566d8066;
mem[2831] = 80'h0010deee97bfbc9cf833;
mem[2832] = 80'h011064b761951bfc167f;
mem[2833] = 80'h00000000000000000000;
mem[2834] = 80'h00000000000000000000;
mem[2835] = 80'h00000000000000000000;
mem[2836] = 80'h10100000010000010010;
mem[2837] = 80'h00109400000208004500;
mem[2838] = 80'h0010002e29f00000fffd;
mem[2839] = 80'h00100f8ac0550102c000;
mem[2840] = 80'h00100001ffabffabffab;
mem[2841] = 80'h00100f3856f97ab5f9a4;
mem[2842] = 80'h001061255a39516ed656;
mem[2843] = 80'h011011ec306406146ca6;
mem[2844] = 80'h00000000000000000000;
mem[2845] = 80'h10100000010000010010;
mem[2846] = 80'h00109400000208004500;
mem[2847] = 80'h0010002e29f10000fffd;
mem[2848] = 80'h00100f89c0550102c000;
mem[2849] = 80'h00100001ffabffabffab;
mem[2850] = 80'h00100e4988d5a2cc3b1b;
mem[2851] = 80'h0010aaf7ddd4a4be9707;
mem[2852] = 80'h01105edb678b9f64e8e0;
mem[2853] = 80'h00000000000000000000;
mem[2854] = 80'h00000000000000000000;
mem[2855] = 80'h00000000000000000000;
mem[2856] = 80'h10100000010000010010;
mem[2857] = 80'h00109400000208004500;
mem[2858] = 80'h0010002e29f20000fffd;
mem[2859] = 80'h00100f88c0550102c000;
mem[2860] = 80'h00100001ffabffabffab;
mem[2861] = 80'h00100ddbeaa0ca467cdb;
mem[2862] = 80'h0010f68055e2bace52f5;
mem[2863] = 80'h01103505313569482cad;
mem[2864] = 80'h00000000000000000000;
mem[2865] = 80'h10100000010000010010;
mem[2866] = 80'h00109400000208004500;
mem[2867] = 80'h0010002e29f30000fffd;
mem[2868] = 80'h00100f87c0550102c000;
mem[2869] = 80'h00100001ffabffabffab;
mem[2870] = 80'h00100caa348c123fbe64;
mem[2871] = 80'h00103d52d20f4f1e2ba4;
mem[2872] = 80'h0110f60e6df2d12be11d;
mem[2873] = 80'h00000000000000000000;
mem[2874] = 80'h00000000000000000000;
mem[2875] = 80'h00000000000000000000;
mem[2876] = 80'h00000000000000000000;
mem[2877] = 80'h10100000010000010010;
mem[2878] = 80'h00109400000208004500;
mem[2879] = 80'h0010002e29f40000fffd;
mem[2880] = 80'h00100f86c0550102c000;
mem[2881] = 80'h00100001ffabffabffab;
mem[2882] = 80'h00100b8ef066c32b31e4;
mem[2883] = 80'h001085bdc36373ff5241;
mem[2884] = 80'h01100190fe08bb4cf688;
mem[2885] = 80'h00000000000000000000;
mem[2886] = 80'h00000000000000000000;
mem[2887] = 80'h00000000000000000000;
mem[2888] = 80'h00000000000000000000;
mem[2889] = 80'h10100000010000010010;
mem[2890] = 80'h00109400000208004500;
mem[2891] = 80'h0010002e29f50000fffd;
mem[2892] = 80'h00100f85c0550102c000;
mem[2893] = 80'h00100001ffabffabffab;
mem[2894] = 80'h00100aff2e4a1b52f35b;
mem[2895] = 80'h00104e6f448e862fdb10;
mem[2896] = 80'h0110d15af26f073edad1;
mem[2897] = 80'h00000000000000000000;
mem[2898] = 80'h00000000000000000000;
mem[2899] = 80'h00000000000000000000;
mem[2900] = 80'h10100000010000010010;
mem[2901] = 80'h00109400000208004500;
mem[2902] = 80'h0010002e29f60000fffd;
mem[2903] = 80'h00100f84c0550102c000;
mem[2904] = 80'h00100001ffabffabffab;
mem[2905] = 80'h0010096d4c3f73d8b49b;
mem[2906] = 80'h00101218ccb8985f50e2;
mem[2907] = 80'h0110944725851eb5d634;
mem[2908] = 80'h00000000000000000000;
mem[2909] = 80'h10100000010000010010;
mem[2910] = 80'h00109400000208004500;
mem[2911] = 80'h0010002e29f70000fffd;
mem[2912] = 80'h00100f83c0550102c000;
mem[2913] = 80'h00100001ffabffabffab;
mem[2914] = 80'h0010081c9213aba17624;
mem[2915] = 80'h0010d9ca4b556d8f4fb3;
mem[2916] = 80'h0110f6c06ae603215f3d;
mem[2917] = 80'h00000000000000000000;
mem[2918] = 80'h00000000000000000000;
mem[2919] = 80'h00000000000000000000;
mem[2920] = 80'h10100000010000010010;
mem[2921] = 80'h00109400000208004500;
mem[2922] = 80'h0010002e29f80000fffd;
mem[2923] = 80'h00100f82c0550102c000;
mem[2924] = 80'h00100001ffabffabffab;
mem[2925] = 80'h00100724c5ead1f1ab9a;
mem[2926] = 80'h001063c6ee60e19dba29;
mem[2927] = 80'h0110c29004e5de32abaf;
mem[2928] = 80'h00000000000000000000;
mem[2929] = 80'h10100000010000010010;
mem[2930] = 80'h00109400000208004500;
mem[2931] = 80'h0010002e29f90000fffd;
mem[2932] = 80'h00100f81c0550102c000;
mem[2933] = 80'h00100001ffabffabffab;
mem[2934] = 80'h001006551bc609886925;
mem[2935] = 80'h0010a814698d144c3a78;
mem[2936] = 80'h01109ff26adeda6cb18a;
mem[2937] = 80'h00000000000000000000;
mem[2938] = 80'h00000000000000000000;
mem[2939] = 80'h00000000000000000000;
mem[2940] = 80'h10100000010000010010;
mem[2941] = 80'h00109400000208004500;
mem[2942] = 80'h0010002e29fa0000fffd;
mem[2943] = 80'h00100f80c0550102c000;
mem[2944] = 80'h00100001ffabffabffab;
mem[2945] = 80'h001005c779b361022ee5;
mem[2946] = 80'h0010f463e1bb0a3c8e8a;
mem[2947] = 80'h0110cf44b272fdbf5c30;
mem[2948] = 80'h00000000000000000000;
mem[2949] = 80'h00000000000000000000;
mem[2950] = 80'h00000000000000000000;
mem[2951] = 80'h10100000010000010010;
mem[2952] = 80'h00109400000208004500;
mem[2953] = 80'h0010002e29fb0000fffd;
mem[2954] = 80'h00100f7fc0550102c000;
mem[2955] = 80'h00100001ffabffabffab;
mem[2956] = 80'h001004b6a79fb97bec5a;
mem[2957] = 80'h00103fb16656ffecc5db;
mem[2958] = 80'h01106fb8d24a02221d28;
mem[2959] = 80'h00000000000000000000;
mem[2960] = 80'h00000000000000000000;
mem[2961] = 80'h00000000000000000000;
mem[2962] = 80'h10100000010000010010;
mem[2963] = 80'h00109400000208004500;
mem[2964] = 80'h0010002e29fc0000fffd;
mem[2965] = 80'h00100f7ec0550102c000;
mem[2966] = 80'h00100001ffabffabffab;
mem[2967] = 80'h001003926375686f63da;
mem[2968] = 80'h0010875e773ac30dfe3e;
mem[2969] = 80'h0110f388194027cb840f;
mem[2970] = 80'h00000000000000000000;
mem[2971] = 80'h10100000010000010010;
mem[2972] = 80'h00109400000208004500;
mem[2973] = 80'h0010002e29fd0000fffd;
mem[2974] = 80'h00100f7dc0550102c000;
mem[2975] = 80'h00100001ffabffabffab;
mem[2976] = 80'h001002e3bd59b016a165;
mem[2977] = 80'h00104c8cf0d736dda16f;
mem[2978] = 80'h01109cc33bd26d66f9f1;
mem[2979] = 80'h00000000000000000000;
mem[2980] = 80'h00000000000000000000;
mem[2981] = 80'h00000000000000000000;
mem[2982] = 80'h00000000000000000000;
mem[2983] = 80'h10100000010000010010;
mem[2984] = 80'h00109400000208004500;
mem[2985] = 80'h0010002e29fe0000fffd;
mem[2986] = 80'h00100f7cc0550102c000;
mem[2987] = 80'h00100001ffabffabffab;
mem[2988] = 80'h00100171df2cd89ce6a5;
mem[2989] = 80'h001010fb78e128ade29d;
mem[2990] = 80'h0110462384d4202fe9b5;
mem[2991] = 80'h00000000000000000000;
mem[2992] = 80'h00000000000000000000;
mem[2993] = 80'h00000000000000000000;
mem[2994] = 80'h10100000010000010010;
mem[2995] = 80'h00109400000208004500;
mem[2996] = 80'h0010002e29ff0000fffd;
mem[2997] = 80'h00100f7bc0550102c000;
mem[2998] = 80'h00100001ffabffabffab;
mem[2999] = 80'h00100000010000e5241a;
mem[3000] = 80'h0010db29ff0cdd7da1cc;
mem[3001] = 80'h01106f761109cdfe3a52;
mem[3002] = 80'h00000000000000000000;
mem[3003] = 80'h10100000010000010010;
mem[3004] = 80'h00109400000208004500;
mem[3005] = 80'h0010002e2a000000fffd;
mem[3006] = 80'h00100f7ac0550102c000;
mem[3007] = 80'h00100001ffabffabffab;
mem[3008] = 80'h0010ff2f4b1bb732658f;
mem[3009] = 80'h00109d9b82578e326003;
mem[3010] = 80'h0110d9a9b11f979030e6;
mem[3011] = 80'h00000000000000000000;
mem[3012] = 80'h00000000000000000000;
mem[3013] = 80'h00000000000000000000;
mem[3014] = 80'h00000000000000000000;
mem[3015] = 80'h10100000010000010010;
mem[3016] = 80'h00109400000208004500;
mem[3017] = 80'h0010002e2a010000fffd;
mem[3018] = 80'h00100f79c0550102c000;
mem[3019] = 80'h00100001ffabffabffab;
mem[3020] = 80'h0010fe5e95376f4ba730;
mem[3021] = 80'h0010564905ba7be26052;
mem[3022] = 80'h0110a8637551711ce532;
mem[3023] = 80'h00000000000000000000;
mem[3024] = 80'h00000000000000000000;
mem[3025] = 80'h00000000000000000000;
mem[3026] = 80'h10100000010000010010;
mem[3027] = 80'h00109400000208004500;
mem[3028] = 80'h0010002e2a020000fffd;
mem[3029] = 80'h00100f78c0550102c000;
mem[3030] = 80'h00100001ffabffabffab;
mem[3031] = 80'h0010fdccf74207c1e0f0;
mem[3032] = 80'h00100a3e8d8c6592e5a0;
mem[3033] = 80'h0110ce7170cedb9359c7;
mem[3034] = 80'h00000000000000000000;
mem[3035] = 80'h10100000010000010010;
mem[3036] = 80'h00109400000208004500;
mem[3037] = 80'h0010002e2a030000fffd;
mem[3038] = 80'h00100f77c0550102c000;
mem[3039] = 80'h00100001ffabffabffab;
mem[3040] = 80'h0010fcbd296edfb8224f;
mem[3041] = 80'h0010c1ec0a6190417df1;
mem[3042] = 80'h011077a985a132c5e1b7;
mem[3043] = 80'h00000000000000000000;
mem[3044] = 80'h00000000000000000000;
mem[3045] = 80'h00000000000000000000;
mem[3046] = 80'h10100000010000010010;
mem[3047] = 80'h00109400000208004500;
mem[3048] = 80'h0010002e2a040000fffd;
mem[3049] = 80'h00100f76c0550102c000;
mem[3050] = 80'h00100001ffabffabffab;
mem[3051] = 80'h0010fb99ed840eacadcf;
mem[3052] = 80'h001079031b0daca00514;
mem[3053] = 80'h0110b3066199b8e5893b;
mem[3054] = 80'h00000000000000000000;
mem[3055] = 80'h10100000010000010010;
mem[3056] = 80'h00109400000208004500;
mem[3057] = 80'h0010002e2a050000fffd;
mem[3058] = 80'h00100f75c0550102c000;
mem[3059] = 80'h00100001ffabffabffab;
mem[3060] = 80'h0010fae833a8d6d56f70;
mem[3061] = 80'h0010b2d19ce059700d45;
mem[3062] = 80'h01104b65895bc8d0c898;
mem[3063] = 80'h00000000000000000000;
mem[3064] = 80'h00000000000000000000;
mem[3065] = 80'h00000000000000000000;
mem[3066] = 80'h00000000000000000000;
mem[3067] = 80'h10100000010000010010;
mem[3068] = 80'h00109400000208004500;
mem[3069] = 80'h0010002e2a060000fffd;
mem[3070] = 80'h00100f74c0550102c000;
mem[3071] = 80'h00100001ffabffabffab;
mem[3072] = 80'h0010f97a51ddbe5f28b0;
mem[3073] = 80'h0010eea614d64700b8b7;
mem[3074] = 80'h011028e2a180800d93f4;
mem[3075] = 80'h00000000000000000000;
mem[3076] = 80'h00000000000000000000;
mem[3077] = 80'h00000000000000000000;
mem[3078] = 80'h10100000010000010010;
mem[3079] = 80'h00109400000208004500;
mem[3080] = 80'h0010002e2a070000fffd;
mem[3081] = 80'h00100f73c0550102c000;
mem[3082] = 80'h00100001ffabffabffab;
mem[3083] = 80'h0010f80b8ff16626ea0f;
mem[3084] = 80'h00102574933bb2d0f9e6;
mem[3085] = 80'h011067d55a8f263f3598;
mem[3086] = 80'h00000000000000000000;
mem[3087] = 80'h00000000000000000000;
mem[3088] = 80'h00000000000000000000;
mem[3089] = 80'h10100000010000010010;
mem[3090] = 80'h00109400000208004500;
mem[3091] = 80'h0010002e2a080000fffd;
mem[3092] = 80'h00100f72c0550102c000;
mem[3093] = 80'h00100001ffabffabffab;
mem[3094] = 80'h0010f733d8081c7637b1;
mem[3095] = 80'h00109f78360e3ec2cd7c;
mem[3096] = 80'h011076e083f5ca46d88b;
mem[3097] = 80'h00000000000000000000;
mem[3098] = 80'h10100000010000010010;
mem[3099] = 80'h00109400000208004500;
mem[3100] = 80'h0010002e2a090000fffd;
mem[3101] = 80'h00100f71c0550102c000;
mem[3102] = 80'h00100001ffabffabffab;
mem[3103] = 80'h0010f6420624c40ff50e;
mem[3104] = 80'h001054aab1e3cb128c2d;
mem[3105] = 80'h011039d7b2d4c5152782;
mem[3106] = 80'h00000000000000000000;
mem[3107] = 80'h00000000000000000000;
mem[3108] = 80'h00000000000000000000;
mem[3109] = 80'h10100000010000010010;
mem[3110] = 80'h00109400000208004500;
mem[3111] = 80'h0010002e2a0a0000fffd;
mem[3112] = 80'h00100f70c0550102c000;
mem[3113] = 80'h00100001ffabffabffab;
mem[3114] = 80'h0010f5d06451ac85b2ce;
mem[3115] = 80'h001008dd39d5d56259df;
mem[3116] = 80'h0110517a831a13ce8ef2;
mem[3117] = 80'h00000000000000000000;
mem[3118] = 80'h10100000010000010010;
mem[3119] = 80'h00109400000208004500;
mem[3120] = 80'h0010002e2a0b0000fffd;
mem[3121] = 80'h00100f6fc0550102c000;
mem[3122] = 80'h00100001ffabffabffab;
mem[3123] = 80'h0010f4a1ba7d74fc7071;
mem[3124] = 80'h0010c30fbe3820b2138e;
mem[3125] = 80'h0110c2b7f3314ebcf541;
mem[3126] = 80'h00000000000000000000;
mem[3127] = 80'h00000000000000000000;
mem[3128] = 80'h00000000000000000000;
mem[3129] = 80'h10100000010000010010;
mem[3130] = 80'h00109400000208004500;
mem[3131] = 80'h0010002e2a0c0000fffd;
mem[3132] = 80'h00100f6ec0550102c000;
mem[3133] = 80'h00100001ffabffabffab;
mem[3134] = 80'h0010f3857e97a5e8fff1;
mem[3135] = 80'h00107be0af541c52a96b;
mem[3136] = 80'h0110411eb5f61f05b784;
mem[3137] = 80'h00000000000000000000;
mem[3138] = 80'h00000000000000000000;
mem[3139] = 80'h00000000000000000000;
mem[3140] = 80'h00000000000000000000;
mem[3141] = 80'h10100000010000010010;
mem[3142] = 80'h00109400000208004500;
mem[3143] = 80'h0010002e2a0d0000fffd;
mem[3144] = 80'h00100f6dc0550102c000;
mem[3145] = 80'h00100001ffabffabffab;
mem[3146] = 80'h0010f2f4a0bb7d913d4e;
mem[3147] = 80'h0010b03228b9e982d03a;
mem[3148] = 80'h011082159cb005aa52be;
mem[3149] = 80'h00000000000000000000;
mem[3150] = 80'h00000000000000000000;
mem[3151] = 80'h00000000000000000000;
mem[3152] = 80'h10100000010000010010;
mem[3153] = 80'h00109400000208004500;
mem[3154] = 80'h0010002e2a0e0000fffd;
mem[3155] = 80'h00100f6cc0550102c000;
mem[3156] = 80'h00100001ffabffabffab;
mem[3157] = 80'h0010f166c2ce151b7a8e;
mem[3158] = 80'h0010ec45a08ff7f254c8;
mem[3159] = 80'h0110d7360b59731294bd;
mem[3160] = 80'h00000000000000000000;
mem[3161] = 80'h00000000000000000000;
mem[3162] = 80'h00000000000000000000;
mem[3163] = 80'h10100000010000010010;
mem[3164] = 80'h00109400000208004500;
mem[3165] = 80'h0010002e2a0f0000fffd;
mem[3166] = 80'h00100f6bc0550102c000;
mem[3167] = 80'h00100001ffabffabffab;
mem[3168] = 80'h0010f0171ce2cd62b831;
mem[3169] = 80'h00102797276202225499;
mem[3170] = 80'h0110a6fc20c063658a20;
mem[3171] = 80'h00000000000000000000;
mem[3172] = 80'h10100000010000010010;
mem[3173] = 80'h00109400000208004500;
mem[3174] = 80'h0010002e2a100000fffd;
mem[3175] = 80'h00100f6ac0550102c000;
mem[3176] = 80'h00100001ffabffabffab;
mem[3177] = 80'h0010ef166d3ce1bac1f3;
mem[3178] = 80'h0010985ceae4efd7bbfc;
mem[3179] = 80'h011073525d9580da0df0;
mem[3180] = 80'h00000000000000000000;
mem[3181] = 80'h00000000000000000000;
mem[3182] = 80'h00000000000000000000;
mem[3183] = 80'h10100000010000010010;
mem[3184] = 80'h00109400000208004500;
mem[3185] = 80'h0010002e2a110000fffd;
mem[3186] = 80'h00100f69c0550102c000;
mem[3187] = 80'h00100001ffabffabffab;
mem[3188] = 80'h0010ee67b31039c3034c;
mem[3189] = 80'h0010538e6d091a0734ad;
mem[3190] = 80'h0110093e08eec02923ff;
mem[3191] = 80'h00000000000000000000;
mem[3192] = 80'h10100000010000010010;
mem[3193] = 80'h00109400000208004500;
mem[3194] = 80'h0010002e2a120000fffd;
mem[3195] = 80'h00100f68c0550102c000;
mem[3196] = 80'h00100001ffabffabffab;
mem[3197] = 80'h0010edf5d1655149448c;
mem[3198] = 80'h00100ff9e53f0477bf5f;
mem[3199] = 80'h01104c23a59b70bd4faf;
mem[3200] = 80'h00000000000000000000;
mem[3201] = 80'h00000000000000000000;
mem[3202] = 80'h00000000000000000000;
mem[3203] = 80'h00000000000000000000;
mem[3204] = 80'h10100000010000010010;
mem[3205] = 80'h00109400000208004500;
mem[3206] = 80'h0010002e2a130000fffd;
mem[3207] = 80'h00100f67c0550102c000;
mem[3208] = 80'h00100001ffabffabffab;
mem[3209] = 80'h0010ec840f4989308633;
mem[3210] = 80'h0010c42b62d2f1a7c40e;
mem[3211] = 80'h0110e94a2ecee2692cd7;
mem[3212] = 80'h00000000000000000000;
mem[3213] = 80'h00000000000000000000;
mem[3214] = 80'h00000000000000000000;
mem[3215] = 80'h10100000010000010010;
mem[3216] = 80'h00109400000208004500;
mem[3217] = 80'h0010002e2a140000fffd;
mem[3218] = 80'h00100f66c0550102c000;
mem[3219] = 80'h00100001ffabffabffab;
mem[3220] = 80'h0010eba0cba3582409b3;
mem[3221] = 80'h00107cc473becd46ffeb;
mem[3222] = 80'h0110757ab3b38a9e35d2;
mem[3223] = 80'h00000000000000000000;
mem[3224] = 80'h00000000000000000000;
mem[3225] = 80'h00000000000000000000;
mem[3226] = 80'h10100000010000010010;
mem[3227] = 80'h00109400000208004500;
mem[3228] = 80'h0010002e2a150000fffd;
mem[3229] = 80'h00100f65c0550102c000;
mem[3230] = 80'h00100001ffabffabffab;
mem[3231] = 80'h0010ead1158f805dcb0c;
mem[3232] = 80'h0010b716f4533896b0ba;
mem[3233] = 80'h01101942063730e148a1;
mem[3234] = 80'h00000000000000000000;
mem[3235] = 80'h10100000010000010010;
mem[3236] = 80'h00109400000208004500;
mem[3237] = 80'h0010002e2a160000fffd;
mem[3238] = 80'h00100f64c0550102c000;
mem[3239] = 80'h00100001ffabffabffab;
mem[3240] = 80'h0010e94377fae8d78ccc;
mem[3241] = 80'h0010eb617c652619e248;
mem[3242] = 80'h01103c837c70584b38ef;
mem[3243] = 80'h00000000000000000000;
mem[3244] = 80'h00000000000000000000;
mem[3245] = 80'h00000000000000000000;
mem[3246] = 80'h10100000010000010010;
mem[3247] = 80'h00109400000208004500;
mem[3248] = 80'h0010002e2a170000fffd;
mem[3249] = 80'h00100f63c0550102c000;
mem[3250] = 80'h00100001ffabffabffab;
mem[3251] = 80'h0010e832a9d630ae4e73;
mem[3252] = 80'h001020b3fb88d3c9a019;
mem[3253] = 80'h011026e737ce8b4980cf;
mem[3254] = 80'h00000000000000000000;
mem[3255] = 80'h00000000000000000000;
mem[3256] = 80'h00000000000000000000;
mem[3257] = 80'h10100000010000010010;
mem[3258] = 80'h00109400000208004500;
mem[3259] = 80'h0010002e2a180000fffd;
mem[3260] = 80'h00100f62c0550102c000;
mem[3261] = 80'h00100001ffabffabffab;
mem[3262] = 80'h0010e70afe2f4afe93cd;
mem[3263] = 80'h00109abf5ebd5fdb1783;
mem[3264] = 80'h01107919520486526921;
mem[3265] = 80'h00000000000000000000;
mem[3266] = 80'h10100000010000010010;
mem[3267] = 80'h00109400000208004500;
mem[3268] = 80'h0010002e2a190000fffd;
mem[3269] = 80'h00100f61c0550102c000;
mem[3270] = 80'h00100001ffabffabffab;
mem[3271] = 80'h0010e67b200392875172;
mem[3272] = 80'h0010516dd950aa0b56d2;
mem[3273] = 80'h0110362eb3bc76ef7d20;
mem[3274] = 80'h00000000000000000000;
mem[3275] = 80'h00000000000000000000;
mem[3276] = 80'h00000000000000000000;
mem[3277] = 80'h00000000000000000000;
mem[3278] = 80'h10100000010000010010;
mem[3279] = 80'h00109400000208004500;
mem[3280] = 80'h0010002e2a1a0000fffd;
mem[3281] = 80'h00100f60c0550102c000;
mem[3282] = 80'h00100001ffabffabffab;
mem[3283] = 80'h0010e5e94276fa0d16b2;
mem[3284] = 80'h00100d1a5166b47be220;
mem[3285] = 80'h011066986b2ae3e59c5c;
mem[3286] = 80'h00000000000000000000;
mem[3287] = 80'h10100000010000010010;
mem[3288] = 80'h00109400000208004500;
mem[3289] = 80'h0010002e2a1b0000fffd;
mem[3290] = 80'h00100f5fc0550102c000;
mem[3291] = 80'h00100001ffabffabffab;
mem[3292] = 80'h0010e4989c5a2274d40d;
mem[3293] = 80'h0010c6c8d68b41ab6a71;
mem[3294] = 80'h01108563b9b5d730d737;
mem[3295] = 80'h00000000000000000000;
mem[3296] = 80'h00000000000000000000;
mem[3297] = 80'h00000000000000000000;
mem[3298] = 80'h00000000000000000000;
mem[3299] = 80'h10100000010000010010;
mem[3300] = 80'h00109400000208004500;
mem[3301] = 80'h0010002e2a1c0000fffd;
mem[3302] = 80'h00100f5ec0550102c000;
mem[3303] = 80'h00100001ffabffabffab;
mem[3304] = 80'h0010e3bc58b0f3605b8d;
mem[3305] = 80'h00107e27c7e77d4a1394;
mem[3306] = 80'h011072fd2ab994001ef6;
mem[3307] = 80'h00000000000000000000;
mem[3308] = 80'h00000000000000000000;
mem[3309] = 80'h00000000000000000000;
mem[3310] = 80'h10100000010000010010;
mem[3311] = 80'h00109400000208004500;
mem[3312] = 80'h0010002e2a1d0000fffd;
mem[3313] = 80'h00100f5dc0550102c000;
mem[3314] = 80'h00100001ffabffabffab;
mem[3315] = 80'h0010e2cd869c2b199932;
mem[3316] = 80'h0010b5f5400a889a0ac5;
mem[3317] = 80'h0110badc8e0dd5914afb;
mem[3318] = 80'h00000000000000000000;
mem[3319] = 80'h10100000010000010010;
mem[3320] = 80'h00109400000208004500;
mem[3321] = 80'h0010002e2a1e0000fffd;
mem[3322] = 80'h00100f5cc0550102c000;
mem[3323] = 80'h00100001ffabffabffab;
mem[3324] = 80'h0010e15fe4e94393def2;
mem[3325] = 80'h0010e982c83c96ea8f37;
mem[3326] = 80'h0110dcce627f1fc8f15f;
mem[3327] = 80'h00000000000000000000;
mem[3328] = 80'h00000000000000000000;
mem[3329] = 80'h00000000000000000000;
mem[3330] = 80'h10100000010000010010;
mem[3331] = 80'h00109400000208004500;
mem[3332] = 80'h0010002e2a1f0000fffd;
mem[3333] = 80'h00100f5bc0550102c000;
mem[3334] = 80'h00100001ffabffabffab;
mem[3335] = 80'h0010e02e3ac59bea1c4d;
mem[3336] = 80'h001022504fd1633b0e66;
mem[3337] = 80'h0110b29d96736b0909cd;
mem[3338] = 80'h00000000000000000000;
mem[3339] = 80'h00000000000000000000;
mem[3340] = 80'h00000000000000000000;
mem[3341] = 80'h10100000010000010010;
mem[3342] = 80'h00109400000208004500;
mem[3343] = 80'h0010002e2a200000fffd;
mem[3344] = 80'h00100f5ac0550102c000;
mem[3345] = 80'h00100001ffabffabffab;
mem[3346] = 80'h0010df5d07551a232d77;
mem[3347] = 80'h0010961553314d00d5fd;
mem[3348] = 80'h011087df3d8ec6de333b;
mem[3349] = 80'h00000000000000000000;
mem[3350] = 80'h10100000010000010010;
mem[3351] = 80'h00109400000208004500;
mem[3352] = 80'h0010002e2a210000fffd;
mem[3353] = 80'h00100f59c0550102c000;
mem[3354] = 80'h00100001ffabffabffab;
mem[3355] = 80'h0010de2cd979c25aefc8;
mem[3356] = 80'h00105dc7d4dcb8d09bac;
mem[3357] = 80'h0110d8d6363d088cde86;
mem[3358] = 80'h00000000000000000000;
mem[3359] = 80'h00000000000000000000;
mem[3360] = 80'h00000000000000000000;
mem[3361] = 80'h00000000000000000000;
mem[3362] = 80'h10100000010000010010;
mem[3363] = 80'h00109400000208004500;
mem[3364] = 80'h0010002e2a220000fffd;
mem[3365] = 80'h00100f58c0550102c000;
mem[3366] = 80'h00100001ffabffabffab;
mem[3367] = 80'h0010ddbebb0caad0a808;
mem[3368] = 80'h001001b05ceaa6a0515e;
mem[3369] = 80'h0110a3361a8b6094ab9f;
mem[3370] = 80'h00000000000000000000;
mem[3371] = 80'h00000000000000000000;
mem[3372] = 80'h00000000000000000000;
mem[3373] = 80'h10100000010000010010;
mem[3374] = 80'h00109400000208004500;
mem[3375] = 80'h0010002e2a230000fffd;
mem[3376] = 80'h00100f57c0550102c000;
mem[3377] = 80'h00100001ffabffabffab;
mem[3378] = 80'h0010dccf652072a96ab7;
mem[3379] = 80'h0010ca62db0753700b0f;
mem[3380] = 80'h01103388a93ce882903d;
mem[3381] = 80'h00000000000000000000;
mem[3382] = 80'h10100000010000010010;
mem[3383] = 80'h00109400000208004500;
mem[3384] = 80'h0010002e2a240000fffd;
mem[3385] = 80'h00100f56c0550102c000;
mem[3386] = 80'h00100001ffabffabffab;
mem[3387] = 80'h0010dbeba1caa3bde537;
mem[3388] = 80'h0010728dca6b6f91beea;
mem[3389] = 80'h0110972ff6ae36348918;
mem[3390] = 80'h00000000000000000000;
mem[3391] = 80'h00000000000000000000;
mem[3392] = 80'h00000000000000000000;
mem[3393] = 80'h10100000010000010010;
mem[3394] = 80'h00109400000208004500;
mem[3395] = 80'h0010002e2a250000fffd;
mem[3396] = 80'h00100f55c0550102c000;
mem[3397] = 80'h00100001ffabffabffab;
mem[3398] = 80'h0010da9a7fe67bc42788;
mem[3399] = 80'h0010b95f4d869a41f8bb;
mem[3400] = 80'h0110418f26bfdba5db55;
mem[3401] = 80'h00000000000000000000;
mem[3402] = 80'h00000000000000000000;
mem[3403] = 80'h00000000000000000000;
mem[3404] = 80'h10100000010000010010;
mem[3405] = 80'h00109400000208004500;
mem[3406] = 80'h0010002e2a260000fffd;
mem[3407] = 80'h00100f54c0550102c000;
mem[3408] = 80'h00100001ffabffabffab;
mem[3409] = 80'h0010d9081d93134e6048;
mem[3410] = 80'h0010e528c5b084314c49;
mem[3411] = 80'h011011390940c801a946;
mem[3412] = 80'h00000000000000000000;
mem[3413] = 80'h00000000000000000000;
mem[3414] = 80'h00000000000000000000;
mem[3415] = 80'h10100000010000010010;
mem[3416] = 80'h00109400000208004500;
mem[3417] = 80'h0010002e2a270000fffd;
mem[3418] = 80'h00100f53c0550102c000;
mem[3419] = 80'h00100001ffabffabffab;
mem[3420] = 80'h0010d879c3bfcb37a2f7;
mem[3421] = 80'h00102efa425d71e14f18;
mem[3422] = 80'h011035a08da53ef626bf;
mem[3423] = 80'h00000000000000000000;
mem[3424] = 80'h10100000010000010010;
mem[3425] = 80'h00109400000208004500;
mem[3426] = 80'h0010002e2a280000fffd;
mem[3427] = 80'h00100f52c0550102c000;
mem[3428] = 80'h00100001ffabffabffab;
mem[3429] = 80'h0010d7419446b1677f49;
mem[3430] = 80'h001094f6e768fdf3b982;
mem[3431] = 80'h011054a3db4ca94f2f6e;
mem[3432] = 80'h00000000000000000000;
mem[3433] = 80'h00000000000000000000;
mem[3434] = 80'h00000000000000000000;
mem[3435] = 80'h00000000000000000000;
mem[3436] = 80'h10100000010000010010;
mem[3437] = 80'h00109400000208004500;
mem[3438] = 80'h0010002e2a290000fffd;
mem[3439] = 80'h00100f51c0550102c000;
mem[3440] = 80'h00100001ffabffabffab;
mem[3441] = 80'h0010d6304a6a691ebdf6;
mem[3442] = 80'h00105f246085082026d3;
mem[3443] = 80'h011074ec54c68f5ce97c;
mem[3444] = 80'h00000000000000000000;
mem[3445] = 80'h10100000010000010010;
mem[3446] = 80'h00109400000208004500;
mem[3447] = 80'h0010002e2a2a0000fffd;
mem[3448] = 80'h00100f50c0550102c000;
mem[3449] = 80'h00100001ffabffabffab;
mem[3450] = 80'h0010d5a2281f0194fa36;
mem[3451] = 80'h00100353e8b31650ad21;
mem[3452] = 80'h011031f12509be18bc2a;
mem[3453] = 80'h00000000000000000000;
mem[3454] = 80'h00000000000000000000;
mem[3455] = 80'h00000000000000000000;
mem[3456] = 80'h00000000000000000000;
mem[3457] = 80'h10100000010000010010;
mem[3458] = 80'h00109400000208004500;
mem[3459] = 80'h0010002e2a2b0000fffd;
mem[3460] = 80'h00100f4fc0550102c000;
mem[3461] = 80'h00100001ffabffabffab;
mem[3462] = 80'h0010d4d3f633d9ed3889;
mem[3463] = 80'h0010c8816f5ee380a670;
mem[3464] = 80'h01109cc1c3ed862eebdc;
mem[3465] = 80'h00000000000000000000;
mem[3466] = 80'h00000000000000000000;
mem[3467] = 80'h00000000000000000000;
mem[3468] = 80'h10100000010000010010;
mem[3469] = 80'h00109400000208004500;
mem[3470] = 80'h0010002e2a2c0000fffd;
mem[3471] = 80'h00100f4ec0550102c000;
mem[3472] = 80'h00100001ffabffabffab;
mem[3473] = 80'h0010d3f732d908f9b709;
mem[3474] = 80'h0010706e7e32df61dc95;
mem[3475] = 80'h01103e0c50877fc74ead;
mem[3476] = 80'h00000000000000000000;
mem[3477] = 80'h10100000010000010010;
mem[3478] = 80'h00109400000208004500;
mem[3479] = 80'h0010002e2a2d0000fffd;
mem[3480] = 80'h00100f4dc0550102c000;
mem[3481] = 80'h00100001ffabffabffab;
mem[3482] = 80'h0010d286ecf5d08075b6;
mem[3483] = 80'h0010bbbcf9df2ab1a2c4;
mem[3484] = 80'h0110649012a98003da77;
mem[3485] = 80'h00000000000000000000;
mem[3486] = 80'h00000000000000000000;
mem[3487] = 80'h00000000000000000000;
mem[3488] = 80'h00000000000000000000;
mem[3489] = 80'h10100000010000010010;
mem[3490] = 80'h00109400000208004500;
mem[3491] = 80'h0010002e2a2e0000fffd;
mem[3492] = 80'h00100f4cc0550102c000;
mem[3493] = 80'h00100001ffabffabffab;
mem[3494] = 80'h0010d1148e80b80a3276;
mem[3495] = 80'h0010e7cb71e934c1e036;
mem[3496] = 80'h01108d41b9faae330e0a;
mem[3497] = 80'h00000000000000000000;
mem[3498] = 80'h10100000010000010010;
mem[3499] = 80'h00109400000208004500;
mem[3500] = 80'h0010002e2a2f0000fffd;
mem[3501] = 80'h00100f4bc0550102c000;
mem[3502] = 80'h00100001ffabffabffab;
mem[3503] = 80'h0010d06550ac6073f0c9;
mem[3504] = 80'h00102c19f604c111a367;
mem[3505] = 80'h0110a4146304fbc05b38;
mem[3506] = 80'h00000000000000000000;
mem[3507] = 80'h00000000000000000000;
mem[3508] = 80'h00000000000000000000;
mem[3509] = 80'h00000000000000000000;
mem[3510] = 80'h10100000010000010010;
mem[3511] = 80'h00109400000208004500;
mem[3512] = 80'h0010002e2a300000fffd;
mem[3513] = 80'h00100f4ac0550102c000;
mem[3514] = 80'h00100001ffabffabffab;
mem[3515] = 80'h0010cf6421724cab890b;
mem[3516] = 80'h001093d23b822ce40f02;
mem[3517] = 80'h011029250512ea0405df;
mem[3518] = 80'h00000000000000000000;
mem[3519] = 80'h00000000000000000000;
mem[3520] = 80'h00000000000000000000;
mem[3521] = 80'h10100000010000010010;
mem[3522] = 80'h00109400000208004500;
mem[3523] = 80'h0010002e2a310000fffd;
mem[3524] = 80'h00100f49c0550102c000;
mem[3525] = 80'h00100001ffabffabffab;
mem[3526] = 80'h0010ce15ff5e94d24bb4;
mem[3527] = 80'h00105800bc6fd9344e53;
mem[3528] = 80'h01106612aff99a2ffe3f;
mem[3529] = 80'h00000000000000000000;
mem[3530] = 80'h10100000010000010010;
mem[3531] = 80'h00109400000208004500;
mem[3532] = 80'h0010002e2a320000fffd;
mem[3533] = 80'h00100f48c0550102c000;
mem[3534] = 80'h00100001ffabffabffab;
mem[3535] = 80'h0010cd879d2bfc580c74;
mem[3536] = 80'h001004773459c7450ba1;
mem[3537] = 80'h011021645f64436a48ad;
mem[3538] = 80'h00000000000000000000;
mem[3539] = 80'h00000000000000000000;
mem[3540] = 80'h00000000000000000000;
mem[3541] = 80'h00000000000000000000;
mem[3542] = 80'h10100000010000010010;
mem[3543] = 80'h00109400000208004500;
mem[3544] = 80'h0010002e2a330000fffd;
mem[3545] = 80'h00100f47c0550102c000;
mem[3546] = 80'h00100001ffabffabffab;
mem[3547] = 80'h0010ccf643072421cecb;
mem[3548] = 80'h0010cfa5b3b4329572f0;
mem[3549] = 80'h0110e26ff1c43f7ed9e8;
mem[3550] = 80'h00000000000000000000;
mem[3551] = 80'h00000000000000000000;
mem[3552] = 80'h00000000000000000000;
mem[3553] = 80'h10100000010000010010;
mem[3554] = 80'h00109400000208004500;
mem[3555] = 80'h0010002e2a340000fffd;
mem[3556] = 80'h00100f46c0550102c000;
mem[3557] = 80'h00100001ffabffabffab;
mem[3558] = 80'h0010cbd287edf535414b;
mem[3559] = 80'h0010774aa2d80e740b15;
mem[3560] = 80'h011015f12c212b763c9e;
mem[3561] = 80'h00000000000000000000;
mem[3562] = 80'h10100000010000010010;
mem[3563] = 80'h00109400000208004500;
mem[3564] = 80'h0010002e2a350000fffd;
mem[3565] = 80'h00100f45c0550102c000;
mem[3566] = 80'h00100001ffabffabffab;
mem[3567] = 80'h0010caa359c12d4c83f4;
mem[3568] = 80'h0010bc982535fba40244;
mem[3569] = 80'h0110dea36bff7fb4880c;
mem[3570] = 80'h00000000000000000000;
mem[3571] = 80'h00000000000000000000;
mem[3572] = 80'h00000000000000000000;
mem[3573] = 80'h10100000010000010010;
mem[3574] = 80'h00109400000208004500;
mem[3575] = 80'h0010002e2a360000fffd;
mem[3576] = 80'h00100f44c0550102c000;
mem[3577] = 80'h00100001ffabffabffab;
mem[3578] = 80'h0010c9313bb445c6c434;
mem[3579] = 80'h0010e0efad03e5d497b6;
mem[3580] = 80'h0110bbc229dd5a5608b4;
mem[3581] = 80'h00000000000000000000;
mem[3582] = 80'h00000000000000000000;
mem[3583] = 80'h00000000000000000000;
mem[3584] = 80'h10100000010000010010;
mem[3585] = 80'h00109400000208004500;
mem[3586] = 80'h0010002e2a370000fffd;
mem[3587] = 80'h00100f43c0550102c000;
mem[3588] = 80'h00100001ffabffabffab;
mem[3589] = 80'h0010c840e5989dbf068b;
mem[3590] = 80'h00102b3d2aee100415e7;
mem[3591] = 80'h0110b7f279d2928ccf8e;
mem[3592] = 80'h00000000000000000000;
mem[3593] = 80'h00000000000000000000;
mem[3594] = 80'h00000000000000000000;
mem[3595] = 80'h10100000010000010010;
mem[3596] = 80'h00109400000208004500;
mem[3597] = 80'h0010002e2a380000fffd;
mem[3598] = 80'h00100f42c0550102c000;
mem[3599] = 80'h00100001ffabffabffab;
mem[3600] = 80'h0010c778b261e7efdb35;
mem[3601] = 80'h001091318fdb9c16e27d;
mem[3602] = 80'h0110e5c03d9d4648ec14;
mem[3603] = 80'h00000000000000000000;
mem[3604] = 80'h10100000010000010010;
mem[3605] = 80'h00109400000208004500;
mem[3606] = 80'h0010002e2a390000fffd;
mem[3607] = 80'h00100f41c0550102c000;
mem[3608] = 80'h00100001ffabffabffab;
mem[3609] = 80'h0010c6096c4d3f96198a;
mem[3610] = 80'h00105ae3083669c69c2c;
mem[3611] = 80'h0110bf5c4c1f4a0673e5;
mem[3612] = 80'h00000000000000000000;
mem[3613] = 80'h00000000000000000000;
mem[3614] = 80'h00000000000000000000;
mem[3615] = 80'h10100000010000010010;
mem[3616] = 80'h00109400000208004500;
mem[3617] = 80'h0010002e2a3a0000fffd;
mem[3618] = 80'h00100f40c0550102c000;
mem[3619] = 80'h00100001ffabffabffab;
mem[3620] = 80'h0010c59b0e38571c5e4a;
mem[3621] = 80'h00100694800077b655de;
mem[3622] = 80'h011091ef90acc7166d8c;
mem[3623] = 80'h00000000000000000000;
mem[3624] = 80'h00000000000000000000;
mem[3625] = 80'h00000000000000000000;
mem[3626] = 80'h10100000010000010010;
mem[3627] = 80'h00109400000208004500;
mem[3628] = 80'h0010002e2a3b0000fffd;
mem[3629] = 80'h00100f3fc0550102c000;
mem[3630] = 80'h00100001ffabffabffab;
mem[3631] = 80'h0010c4ead0148f659cf5;
mem[3632] = 80'h0010cd4607ed82661c8f;
mem[3633] = 80'h01105771730af2c0a299;
mem[3634] = 80'h00000000000000000000;
mem[3635] = 80'h00000000000000000000;
mem[3636] = 80'h00000000000000000000;
mem[3637] = 80'h10100000010000010010;
mem[3638] = 80'h00109400000208004500;
mem[3639] = 80'h0010002e2a3c0000fffd;
mem[3640] = 80'h00100f3ec0550102c000;
mem[3641] = 80'h00100001ffabffabffab;
mem[3642] = 80'h0010c3ce14fe5e711375;
mem[3643] = 80'h001075a91681be80a76a;
mem[3644] = 80'h011055496ded316b5414;
mem[3645] = 80'h00000000000000000000;
mem[3646] = 80'h10100000010000010010;
mem[3647] = 80'h00109400000208004500;
mem[3648] = 80'h0010002e2a3d0000fffd;
mem[3649] = 80'h00100f3dc0550102c000;
mem[3650] = 80'h00100001ffabffabffab;
mem[3651] = 80'h0010c2bfcad28608d1ca;
mem[3652] = 80'h0010be7b916c4b50f83b;
mem[3653] = 80'h01103a024d2326b9c2ba;
mem[3654] = 80'h00000000000000000000;
mem[3655] = 80'h00000000000000000000;
mem[3656] = 80'h00000000000000000000;
mem[3657] = 80'h00000000000000000000;
mem[3658] = 80'h10100000010000010010;
mem[3659] = 80'h00109400000208004500;
mem[3660] = 80'h0010002e2a3e0000fffd;
mem[3661] = 80'h00100f3cc0550102c000;
mem[3662] = 80'h00100001ffabffabffab;
mem[3663] = 80'h0010c12da8a7ee82960a;
mem[3664] = 80'h0010e20c195a55203bc9;
mem[3665] = 80'h0110fb7a89d15d4b61e2;
mem[3666] = 80'h00000000000000000000;
mem[3667] = 80'h00000000000000000000;
mem[3668] = 80'h00000000000000000000;
mem[3669] = 80'h10100000010000010010;
mem[3670] = 80'h00109400000208004500;
mem[3671] = 80'h0010002e2a3f0000fffd;
mem[3672] = 80'h00100f3bc0550102c000;
mem[3673] = 80'h00100001ffabffabffab;
mem[3674] = 80'h0010c05c768b36fb54b5;
mem[3675] = 80'h001029de9eb7a0f07898;
mem[3676] = 80'h0110d22f891892305e13;
mem[3677] = 80'h00000000000000000000;
mem[3678] = 80'h10100000010000010010;
mem[3679] = 80'h00109400000208004500;
mem[3680] = 80'h0010002e2a400000fffd;
mem[3681] = 80'h00100f3ac0550102c000;
mem[3682] = 80'h00100001ffabffabffab;
mem[3683] = 80'h0010bfcbd386ed10f47f;
mem[3684] = 80'h00108a86209a09578bff;
mem[3685] = 80'h01100869423c1d7c52d3;
mem[3686] = 80'h00000000000000000000;
mem[3687] = 80'h00000000000000000000;
mem[3688] = 80'h00000000000000000000;
mem[3689] = 80'h10100000010000010010;
mem[3690] = 80'h00109400000208004500;
mem[3691] = 80'h0010002e2a410000fffd;
mem[3692] = 80'h00100f39c0550102c000;
mem[3693] = 80'h00100001ffabffabffab;
mem[3694] = 80'h0010beba0daa356936c0;
mem[3695] = 80'h00104154a777fc8705ae;
mem[3696] = 80'h011041349b3b406e921e;
mem[3697] = 80'h00000000000000000000;
mem[3698] = 80'h00000000000000000000;
mem[3699] = 80'h00000000000000000000;
mem[3700] = 80'h10100000010000010010;
mem[3701] = 80'h00109400000208004500;
mem[3702] = 80'h0010002e2a420000fffd;
mem[3703] = 80'h00100f38c0550102c000;
mem[3704] = 80'h00100001ffabffabffab;
mem[3705] = 80'h0010bd286fdf5de37100;
mem[3706] = 80'h00101d232f41e2f78f5c;
mem[3707] = 80'h011037180e43fb31bb2b;
mem[3708] = 80'h00000000000000000000;
mem[3709] = 80'h00000000000000000000;
mem[3710] = 80'h00000000000000000000;
mem[3711] = 80'h10100000010000010010;
mem[3712] = 80'h00109400000208004500;
mem[3713] = 80'h0010002e2a430000fffd;
mem[3714] = 80'h00100f37c0550102c000;
mem[3715] = 80'h00100001ffabffabffab;
mem[3716] = 80'h0010bc59b1f3859ab3bf;
mem[3717] = 80'h0010d6f1a8ac1727940d;
mem[3718] = 80'h0110995b942929a0485c;
mem[3719] = 80'h00000000000000000000;
mem[3720] = 80'h10100000010000010010;
mem[3721] = 80'h00109400000208004500;
mem[3722] = 80'h0010002e2a440000fffd;
mem[3723] = 80'h00100f36c0550102c000;
mem[3724] = 80'h00100001ffabffabffab;
mem[3725] = 80'h0010bb7d7519548e3c3f;
mem[3726] = 80'h00106e1eb9c02bc6efe8;
mem[3727] = 80'h011008a7f26598d2409a;
mem[3728] = 80'h00000000000000000000;
mem[3729] = 80'h00000000000000000000;
mem[3730] = 80'h00000000000000000000;
mem[3731] = 80'h10100000010000010010;
mem[3732] = 80'h00109400000208004500;
mem[3733] = 80'h0010002e2a450000fffd;
mem[3734] = 80'h00100f35c0550102c000;
mem[3735] = 80'h00100001ffabffabffab;
mem[3736] = 80'h0010ba0cab358cf7fe80;
mem[3737] = 80'h0010a5cc3e2dde1760b9;
mem[3738] = 80'h011045fba67efd5f272e;
mem[3739] = 80'h00000000000000000000;
mem[3740] = 80'h00000000000000000000;
mem[3741] = 80'h00000000000000000000;
mem[3742] = 80'h10100000010000010010;
mem[3743] = 80'h00109400000208004500;
mem[3744] = 80'h0010002e2a460000fffd;
mem[3745] = 80'h00100f34c0550102c000;
mem[3746] = 80'h00100001ffabffabffab;
mem[3747] = 80'h0010b99ec940e47db940;
mem[3748] = 80'h0010f9bbb61bc067d34b;
mem[3749] = 80'h01108cda0efc00c83242;
mem[3750] = 80'h00000000000000000000;
mem[3751] = 80'h00000000000000000000;
mem[3752] = 80'h00000000000000000000;
mem[3753] = 80'h10100000010000010010;
mem[3754] = 80'h00109400000208004500;
mem[3755] = 80'h0010002e2a470000fffd;
mem[3756] = 80'h00100f33c0550102c000;
mem[3757] = 80'h00100001ffabffabffab;
mem[3758] = 80'h0010b8ef176c3c047bff;
mem[3759] = 80'h0010326931f635b7901a;
mem[3760] = 80'h0110a58fa7df09bf178c;
mem[3761] = 80'h00000000000000000000;
mem[3762] = 80'h10100000010000010010;
mem[3763] = 80'h00109400000208004500;
mem[3764] = 80'h0010002e2a480000fffd;
mem[3765] = 80'h00100f32c0550102c000;
mem[3766] = 80'h00100001ffabffabffab;
mem[3767] = 80'h0010b7d740954654a641;
mem[3768] = 80'h0010886594c3b9a52680;
mem[3769] = 80'h0110c940546ddb7b5017;
mem[3770] = 80'h00000000000000000000;
mem[3771] = 80'h00000000000000000000;
mem[3772] = 80'h00000000000000000000;
mem[3773] = 80'h00000000000000000000;
mem[3774] = 80'h10100000010000010010;
mem[3775] = 80'h00109400000208004500;
mem[3776] = 80'h0010002e2a490000fffd;
mem[3777] = 80'h00100f31c0550102c000;
mem[3778] = 80'h00100001ffabffabffab;
mem[3779] = 80'h0010b6a69eb99e2d64fe;
mem[3780] = 80'h001043b7132e4c7567d1;
mem[3781] = 80'h0110867715d04d8e29c8;
mem[3782] = 80'h00000000000000000000;
mem[3783] = 80'h00000000000000000000;
mem[3784] = 80'h00000000000000000000;
mem[3785] = 80'h10100000010000010010;
mem[3786] = 80'h00109400000208004500;
mem[3787] = 80'h0010002e2a4a0000fffd;
mem[3788] = 80'h00100f30c0550102c000;
mem[3789] = 80'h00100001ffabffabffab;
mem[3790] = 80'h0010b534fcccf6a7233e;
mem[3791] = 80'h00101fc09b1852053223;
mem[3792] = 80'h0110f542ffd34cda3155;
mem[3793] = 80'h00000000000000000000;
mem[3794] = 80'h10100000010000010010;
mem[3795] = 80'h00109400000208004500;
mem[3796] = 80'h0010002e2a4b0000fffd;
mem[3797] = 80'h00100f2fc0550102c000;
mem[3798] = 80'h00100001ffabffabffab;
mem[3799] = 80'h0010b44522e02edee181;
mem[3800] = 80'h0010d4121cf5a7d57872;
mem[3801] = 80'h0110668fa09a0890ea57;
mem[3802] = 80'h00000000000000000000;
mem[3803] = 80'h00000000000000000000;
mem[3804] = 80'h00000000000000000000;
mem[3805] = 80'h10100000010000010010;
mem[3806] = 80'h00109400000208004500;
mem[3807] = 80'h0010002e2a4c0000fffd;
mem[3808] = 80'h00100f2ec0550102c000;
mem[3809] = 80'h00100001ffabffabffab;
mem[3810] = 80'h0010b361e60affca6e01;
mem[3811] = 80'h00106cfd0d999b344297;
mem[3812] = 80'h0110c98ed6d58a17c52b;
mem[3813] = 80'h00000000000000000000;
mem[3814] = 80'h00000000000000000000;
mem[3815] = 80'h00000000000000000000;
mem[3816] = 80'h10100000010000010010;
mem[3817] = 80'h00109400000208004500;
mem[3818] = 80'h0010002e2a4d0000fffd;
mem[3819] = 80'h00100f2dc0550102c000;
mem[3820] = 80'h00100001ffabffabffab;
mem[3821] = 80'h0010b210382627b3acbe;
mem[3822] = 80'h0010a72f8a746ee43cc6;
mem[3823] = 80'h01109312d0f57374fc82;
mem[3824] = 80'h00000000000000000000;
mem[3825] = 80'h00000000000000000000;
mem[3826] = 80'h00000000000000000000;
mem[3827] = 80'h10100000010000010010;
mem[3828] = 80'h00109400000208004500;
mem[3829] = 80'h0010002e2a4e0000fffd;
mem[3830] = 80'h00100f2cc0550102c000;
mem[3831] = 80'h00100001ffabffabffab;
mem[3832] = 80'h0010b1825a534f39eb7e;
mem[3833] = 80'h0010fb5802427094bd34;
mem[3834] = 80'h011039c45449950e13c6;
mem[3835] = 80'h00000000000000000000;
mem[3836] = 80'h10100000010000010010;
mem[3837] = 80'h00109400000208004500;
mem[3838] = 80'h0010002e2a4f0000fffd;
mem[3839] = 80'h00100f2bc0550102c000;
mem[3840] = 80'h00100001ffabffabffab;
mem[3841] = 80'h0010b0f3847f974029c1;
mem[3842] = 80'h0010308a85af85473c65;
mem[3843] = 80'h011039f757ade88876a5;
mem[3844] = 80'h00000000000000000000;
mem[3845] = 80'h00000000000000000000;
mem[3846] = 80'h00000000000000000000;
mem[3847] = 80'h10100000010000010010;
mem[3848] = 80'h00109400000208004500;
mem[3849] = 80'h0010002e2a500000fffd;
mem[3850] = 80'h00100f2ac0550102c000;
mem[3851] = 80'h00100001ffabffabffab;
mem[3852] = 80'h0010aff2f5a1bb985003;
mem[3853] = 80'h00108f41482968b2d600;
mem[3854] = 80'h011013ac25051c83a20c;
mem[3855] = 80'h00000000000000000000;
mem[3856] = 80'h00000000000000000000;
mem[3857] = 80'h00000000000000000000;
mem[3858] = 80'h10100000010000010010;
mem[3859] = 80'h00109400000208004500;
mem[3860] = 80'h0010002e2a510000fffd;
mem[3861] = 80'h00100f29c0550102c000;
mem[3862] = 80'h00100001ffabffabffab;
mem[3863] = 80'h0010ae832b8d63e192bc;
mem[3864] = 80'h00104493cfc49d62df51;
mem[3865] = 80'h0110d8fec54525d5e768;
mem[3866] = 80'h00000000000000000000;
mem[3867] = 80'h00000000000000000000;
mem[3868] = 80'h00000000000000000000;
mem[3869] = 80'h10100000010000010010;
mem[3870] = 80'h00109400000208004500;
mem[3871] = 80'h0010002e2a520000fffd;
mem[3872] = 80'h00100f28c0550102c000;
mem[3873] = 80'h00100001ffabffabffab;
mem[3874] = 80'h0010ad1149f80b6bd57c;
mem[3875] = 80'h001018e447f2831256a3;
mem[3876] = 80'h0110fb81f1ff7db9058b;
mem[3877] = 80'h00000000000000000000;
mem[3878] = 80'h10100000010000010010;
mem[3879] = 80'h00109400000208004500;
mem[3880] = 80'h0010002e2a530000fffd;
mem[3881] = 80'h00100f27c0550102c000;
mem[3882] = 80'h00100001ffabffabffab;
mem[3883] = 80'h0010ac6097d4d31217c3;
mem[3884] = 80'h0010d336c01f76c22ef2;
mem[3885] = 80'h01100bbb8c2e3a71e84f;
mem[3886] = 80'h00000000000000000000;
mem[3887] = 80'h00000000000000000000;
mem[3888] = 80'h00000000000000000000;
mem[3889] = 80'h00000000000000000000;
mem[3890] = 80'h10100000010000010010;
mem[3891] = 80'h00109400000208004500;
mem[3892] = 80'h0010002e2a540000fffd;
mem[3893] = 80'h00100f26c0550102c000;
mem[3894] = 80'h00100001ffabffabffab;
mem[3895] = 80'h0010ab44533e02069843;
mem[3896] = 80'h00106bd9d1734a239417;
mem[3897] = 80'h0110bf228c881a5fdcf9;
mem[3898] = 80'h00000000000000000000;
mem[3899] = 80'h00000000000000000000;
mem[3900] = 80'h00000000000000000000;
mem[3901] = 80'h10100000010000010010;
mem[3902] = 80'h00109400000208004500;
mem[3903] = 80'h0010002e2a550000fffd;
mem[3904] = 80'h00100f25c0550102c000;
mem[3905] = 80'h00100001ffabffabffab;
mem[3906] = 80'h0010aa358d12da7f5afc;
mem[3907] = 80'h0010a00b569ebff3db46;
mem[3908] = 80'h0110d31a2e3c9a94fba9;
mem[3909] = 80'h00000000000000000000;
mem[3910] = 80'h10100000010000010010;
mem[3911] = 80'h00109400000208004500;
mem[3912] = 80'h0010002e2a560000fffd;
mem[3913] = 80'h00100f24c0550102c000;
mem[3914] = 80'h00100001ffabffabffab;
mem[3915] = 80'h0010a9a7ef67b2f51d3c;
mem[3916] = 80'h0010fc7cdea8a18309b4;
mem[3917] = 80'h01102220ee40f37d8bd4;
mem[3918] = 80'h00000000000000000000;
mem[3919] = 80'h00000000000000000000;
mem[3920] = 80'h00000000000000000000;
mem[3921] = 80'h10100000010000010010;
mem[3922] = 80'h00109400000208004500;
mem[3923] = 80'h0010002e2a570000fffd;
mem[3924] = 80'h00100f23c0550102c000;
mem[3925] = 80'h00100001ffabffabffab;
mem[3926] = 80'h0010a8d6314b6a8cdf83;
mem[3927] = 80'h001037ae594554534be5;
mem[3928] = 80'h01103844725daade9575;
mem[3929] = 80'h00000000000000000000;
mem[3930] = 80'h10100000010000010010;
mem[3931] = 80'h00109400000208004500;
mem[3932] = 80'h0010002e2a580000fffd;
mem[3933] = 80'h00100f22c0550102c000;
mem[3934] = 80'h00100001ffabffabffab;
mem[3935] = 80'h0010a7ee66b210dc023d;
mem[3936] = 80'h00108da2fc70d8407c7f;
mem[3937] = 80'h01104b12b45f3d63a10e;
mem[3938] = 80'h00000000000000000000;
mem[3939] = 80'h00000000000000000000;
mem[3940] = 80'h00000000000000000000;
mem[3941] = 80'h00000000000000000000;
mem[3942] = 80'h10100000010000010010;
mem[3943] = 80'h00109400000208004500;
mem[3944] = 80'h0010002e2a590000fffd;
mem[3945] = 80'h00100f21c0550102c000;
mem[3946] = 80'h00100001ffabffabffab;
mem[3947] = 80'h0010a69fb89ec8a5c082;
mem[3948] = 80'h001046707b9d2d90032e;
mem[3949] = 80'h011022bf020e9be43468;
mem[3950] = 80'h00000000000000000000;
mem[3951] = 80'h00000000000000000000;
mem[3952] = 80'h00000000000000000000;
mem[3953] = 80'h10100000010000010010;
mem[3954] = 80'h00109400000208004500;
mem[3955] = 80'h0010002e2a5a0000fffd;
mem[3956] = 80'h00100f20c0550102c000;
mem[3957] = 80'h00100001ffabffabffab;
mem[3958] = 80'h0010a50ddaeba02f8742;
mem[3959] = 80'h00101a07f3ab33e088dc;
mem[3960] = 80'h011067a2268291197816;
mem[3961] = 80'h00000000000000000000;
mem[3962] = 80'h00000000000000000000;
mem[3963] = 80'h00000000000000000000;
mem[3964] = 80'h10100000010000010010;
mem[3965] = 80'h00109400000208004500;
mem[3966] = 80'h0010002e2a5b0000fffd;
mem[3967] = 80'h00100f1fc0550102c000;
mem[3968] = 80'h00100001ffabffabffab;
mem[3969] = 80'h0010a47c04c7785645fd;
mem[3970] = 80'h0010d1d57446c630838d;
mem[3971] = 80'h0110ca923dfb36d77750;
mem[3972] = 80'h00000000000000000000;
mem[3973] = 80'h10100000010000010010;
mem[3974] = 80'h00109400000208004500;
mem[3975] = 80'h0010002e2a5c0000fffd;
mem[3976] = 80'h00100f1ec0550102c000;
mem[3977] = 80'h00100001ffabffabffab;
mem[3978] = 80'h0010a358c02da942ca7d;
mem[3979] = 80'h0010693a652afad1f868;
mem[3980] = 80'h01105b6e0bab9ca4c538;
mem[3981] = 80'h00000000000000000000;
mem[3982] = 80'h00000000000000000000;
mem[3983] = 80'h00000000000000000000;
mem[3984] = 80'h10100000010000010010;
mem[3985] = 80'h00109400000208004500;
mem[3986] = 80'h0010002e2a5d0000fffd;
mem[3987] = 80'h00100f1dc0550102c000;
mem[3988] = 80'h00100001ffabffabffab;
mem[3989] = 80'h0010a2291e01713b08c2;
mem[3990] = 80'h0010a2e8e2c70f016739;
mem[3991] = 80'h01102271a77b340c45f4;
mem[3992] = 80'h00000000000000000000;
mem[3993] = 80'h10100000010000010010;
mem[3994] = 80'h00109400000208004500;
mem[3995] = 80'h0010002e2a5e0000fffd;
mem[3996] = 80'h00100f1cc0550102c000;
mem[3997] = 80'h00100001ffabffabffab;
mem[3998] = 80'h0010a1bb7c7419b14f02;
mem[3999] = 80'h0010fe9f6af11171e7cb;
mem[4000] = 80'h0110bb965ab71cce3912;
mem[4001] = 80'h00000000000000000000;
mem[4002] = 80'h00000000000000000000;
mem[4003] = 80'h00000000000000000000;
mem[4004] = 80'h00000000000000000000;
mem[4005] = 80'h10100000010000010010;
mem[4006] = 80'h00109400000208004500;
mem[4007] = 80'h0010002e2a5f0000fffd;
mem[4008] = 80'h00100f1bc0550102c000;
mem[4009] = 80'h00100001ffabffabffab;
mem[4010] = 80'h0010a0caa258c1c88dbd;
mem[4011] = 80'h0010354ded1ce4a1e79a;
mem[4012] = 80'h0110ca5cb45210a71960;
mem[4013] = 80'h00000000000000000000;
mem[4014] = 80'h00000000000000000000;
mem[4015] = 80'h00000000000000000000;
mem[4016] = 80'h00000000000000000000;
mem[4017] = 80'h10100000010000010010;
mem[4018] = 80'h00109400000208004500;
mem[4019] = 80'h0010002e2a600000fffd;
mem[4020] = 80'h00100f1ac0550102c000;
mem[4021] = 80'h00100001ffabffabffab;
mem[4022] = 80'h00109fb99fc84001bc87;
mem[4023] = 80'h00108108f1fcca9a3e01;
mem[4024] = 80'h0110997caed64630f25a;
mem[4025] = 80'h00000000000000000000;
mem[4026] = 80'h00000000000000000000;
mem[4027] = 80'h00000000000000000000;
mem[4028] = 80'h10100000010000010010;
mem[4029] = 80'h00109400000208004500;
mem[4030] = 80'h0010002e2a610000fffd;
mem[4031] = 80'h00100f19c0550102c000;
mem[4032] = 80'h00100001ffabffabffab;
mem[4033] = 80'h00109ec841e498787e38;
mem[4034] = 80'h00104ada76113f4a7050;
mem[4035] = 80'h0110c675d1a5ca1c2837;
mem[4036] = 80'h00000000000000000000;
mem[4037] = 80'h10100000010000010010;
mem[4038] = 80'h00109400000208004500;
mem[4039] = 80'h0010002e2a620000fffd;
mem[4040] = 80'h00100f18c0550102c000;
mem[4041] = 80'h00100001ffabffabffab;
mem[4042] = 80'h00109d5a2391f0f239f8;
mem[4043] = 80'h001016adfe2721353aa2;
mem[4044] = 80'h01108a3c1940c2f080b5;
mem[4045] = 80'h00000000000000000000;
mem[4046] = 80'h00000000000000000000;
mem[4047] = 80'h00000000000000000000;
mem[4048] = 80'h10100000010000010010;
mem[4049] = 80'h00109400000208004500;
mem[4050] = 80'h0010002e2a630000fffd;
mem[4051] = 80'h00100f17c0550102c000;
mem[4052] = 80'h00100001ffabffabffab;
mem[4053] = 80'h00109c2bfdbd288bfb47;
mem[4054] = 80'h0010dd7f79cad4e560f3;
mem[4055] = 80'h01101a829a9dff589a65;
mem[4056] = 80'h00000000000000000000;
mem[4057] = 80'h10100000010000010010;
mem[4058] = 80'h00109400000208004500;
mem[4059] = 80'h0010002e2a640000fffd;
mem[4060] = 80'h00100f16c0550102c000;
mem[4061] = 80'h00100001ffabffabffab;
mem[4062] = 80'h00109b0f3957f99f74c7;
mem[4063] = 80'h0010659068a6e8045516;
mem[4064] = 80'h0110a5bd0c225df3cc75;
mem[4065] = 80'h00000000000000000000;
mem[4066] = 80'h00000000000000000000;
mem[4067] = 80'h00000000000000000000;
mem[4068] = 80'h10100000010000010010;
mem[4069] = 80'h00109400000208004500;
mem[4070] = 80'h0010002e2a650000fffd;
mem[4071] = 80'h00100f15c0550102c000;
mem[4072] = 80'h00100001ffabffabffab;
mem[4073] = 80'h00109a7ee77b21e6b678;
mem[4074] = 80'h0010ae42ef4b1dd41447;
mem[4075] = 80'h0110ea8aeb71dbd25a15;
mem[4076] = 80'h00000000000000000000;
mem[4077] = 80'h00000000000000000000;
mem[4078] = 80'h00000000000000000000;
mem[4079] = 80'h10100000010000010010;
mem[4080] = 80'h00109400000208004500;
mem[4081] = 80'h0010002e2a660000fffd;
mem[4082] = 80'h00100f14c0550102c000;
mem[4083] = 80'h00100001ffabffabffab;
mem[4084] = 80'h001099ec850e496cf1b8;
mem[4085] = 80'h0010f235677d03a4a5b5;
mem[4086] = 80'h011045c95d096177b0e8;
mem[4087] = 80'h00000000000000000000;
mem[4088] = 80'h00000000000000000000;
mem[4089] = 80'h00000000000000000000;
mem[4090] = 80'h10100000010000010010;
mem[4091] = 80'h00109400000208004500;
mem[4092] = 80'h0010002e2a670000fffd;
mem[4093] = 80'h00100f13c0550102c000;
mem[4094] = 80'h00100001ffabffabffab;
mem[4095] = 80'h0010989d5b2291153307;
mem[4096] = 80'h001039e7e090f67424e4;
mem[4097] = 80'h01101caaf5a7b5487ebb;
mem[4098] = 80'h00000000000000000000;
mem[4099] = 80'h10100000010000010010;
mem[4100] = 80'h00109400000208004500;
mem[4101] = 80'h0010002e2a680000fffd;
mem[4102] = 80'h00100f12c0550102c000;
mem[4103] = 80'h00100001ffabffabffab;
mem[4104] = 80'h001097a50cdbeb45eeb9;
mem[4105] = 80'h001083eb45a57a66d47e;
mem[4106] = 80'h0110d70f91f9d2b878fb;
mem[4107] = 80'h00000000000000000000;
mem[4108] = 80'h00000000000000000000;
mem[4109] = 80'h00000000000000000000;
mem[4110] = 80'h10100000010000010010;
mem[4111] = 80'h00109400000208004500;
mem[4112] = 80'h0010002e2a690000fffd;
mem[4113] = 80'h00100f11c0550102c000;
mem[4114] = 80'h00100001ffabffabffab;
mem[4115] = 80'h001096d4d2f7333c2c06;
mem[4116] = 80'h00104839c2488fb6cc2f;
mem[4117] = 80'h01102c1fa469547d1eae;
mem[4118] = 80'h00000000000000000000;
mem[4119] = 80'h00000000000000000000;
mem[4120] = 80'h00000000000000000000;
mem[4121] = 80'h10100000010000010010;
mem[4122] = 80'h00109400000208004500;
mem[4123] = 80'h0010002e2a6a0000fffd;
mem[4124] = 80'h00100f10c0550102c000;
mem[4125] = 80'h00100001ffabffabffab;
mem[4126] = 80'h00109546b0825bb66bc6;
mem[4127] = 80'h0010144e4a7e91c644dd;
mem[4128] = 80'h01103c5180f850f1e9a7;
mem[4129] = 80'h00000000000000000000;
mem[4130] = 80'h00000000000000000000;
mem[4131] = 80'h00000000000000000000;
mem[4132] = 80'h10100000010000010010;
mem[4133] = 80'h00109400000208004500;
mem[4134] = 80'h0010002e2a6b0000fffd;
mem[4135] = 80'h00100f0fc0550102c000;
mem[4136] = 80'h00100001ffabffabffab;
mem[4137] = 80'h001094376eae83cfa979;
mem[4138] = 80'h0010df9ccd936417cc8c;
mem[4139] = 80'h0110e89a096164a39a0c;
mem[4140] = 80'h00000000000000000000;
mem[4141] = 80'h00000000000000000000;
mem[4142] = 80'h00000000000000000000;
mem[4143] = 80'h00000000000000000000;
mem[4144] = 80'h10100000010000010010;
mem[4145] = 80'h00109400000208004500;
mem[4146] = 80'h0010002e2a6c0000fffd;
mem[4147] = 80'h00100f0ec0550102c000;
mem[4148] = 80'h00100001ffabffabffab;
mem[4149] = 80'h00109313aa4452db26f9;
mem[4150] = 80'h00106773dcff58f6b769;
mem[4151] = 80'h011079667a9954402b31;
mem[4152] = 80'h00000000000000000000;
mem[4153] = 80'h10100000010000010010;
mem[4154] = 80'h00109400000208004500;
mem[4155] = 80'h0010002e2a6d0000fffd;
mem[4156] = 80'h00100f0dc0550102c000;
mem[4157] = 80'h00100001ffabffabffab;
mem[4158] = 80'h0010926274688aa2e446;
mem[4159] = 80'h0010aca15b12ad26c938;
mem[4160] = 80'h011023fae83d8a2bea67;
mem[4161] = 80'h00000000000000000000;
mem[4162] = 80'h00000000000000000000;
mem[4163] = 80'h00000000000000000000;
mem[4164] = 80'h10100000010000010010;
mem[4165] = 80'h00109400000208004500;
mem[4166] = 80'h0010002e2a6e0000fffd;
mem[4167] = 80'h00100f0cc0550102c000;
mem[4168] = 80'h00100001ffabffabffab;
mem[4169] = 80'h001091f0161de228a386;
mem[4170] = 80'h0010f0d6d324b3560bca;
mem[4171] = 80'h0110d1b37d7298715225;
mem[4172] = 80'h00000000000000000000;
mem[4173] = 80'h10100000010000010010;
mem[4174] = 80'h00109400000208004500;
mem[4175] = 80'h0010002e2a6f0000fffd;
mem[4176] = 80'h00100f0bc0550102c000;
mem[4177] = 80'h00100001ffabffabffab;
mem[4178] = 80'h00109081c8313a516139;
mem[4179] = 80'h00103b0454c94686489b;
mem[4180] = 80'h0110f8e6f3eb66ee061a;
mem[4181] = 80'h00000000000000000000;
mem[4182] = 80'h00000000000000000000;
mem[4183] = 80'h00000000000000000000;
mem[4184] = 80'h10100000010000010010;
mem[4185] = 80'h00109400000208004500;
mem[4186] = 80'h0010002e2a700000fffd;
mem[4187] = 80'h00100f0ac0550102c000;
mem[4188] = 80'h00100001ffabffabffab;
mem[4189] = 80'h00108f80b9ef168918fb;
mem[4190] = 80'h001084cf994fab7364fe;
mem[4191] = 80'h01106e4fea2a3725e027;
mem[4192] = 80'h00000000000000000000;
mem[4193] = 80'h10100000010000010010;
mem[4194] = 80'h00109400000208004500;
mem[4195] = 80'h0010002e2a710000fffd;
mem[4196] = 80'h00100f09c0550102c000;
mem[4197] = 80'h00100001ffabffabffab;
mem[4198] = 80'h00108ef167c3cef0da44;
mem[4199] = 80'h00104f1d1ea25ea32baf;
mem[4200] = 80'h01100277658c10c554a4;
mem[4201] = 80'h00000000000000000000;
mem[4202] = 80'h00000000000000000000;
mem[4203] = 80'h00000000000000000000;
mem[4204] = 80'h00000000000000000000;
mem[4205] = 80'h10100000010000010010;
mem[4206] = 80'h00109400000208004500;
mem[4207] = 80'h0010002e2a720000fffd;
mem[4208] = 80'h00100f08c0550102c000;
mem[4209] = 80'h00100001ffabffabffab;
mem[4210] = 80'h00108d6305b6a67a9d84;
mem[4211] = 80'h0010136a969440d3e05d;
mem[4212] = 80'h01104aa61311ab9aa25d;
mem[4213] = 80'h00000000000000000000;
mem[4214] = 80'h00000000000000000000;
mem[4215] = 80'h00000000000000000000;
mem[4216] = 80'h10100000010000010010;
mem[4217] = 80'h00109400000208004500;
mem[4218] = 80'h0010002e2a730000fffd;
mem[4219] = 80'h00100f07c0550102c000;
mem[4220] = 80'h00100001ffabffabffab;
mem[4221] = 80'h00108c12db9a7e035f3b;
mem[4222] = 80'h0010d8b81179b5039b0c;
mem[4223] = 80'h0110efcf91016f40b5f2;
mem[4224] = 80'h00000000000000000000;
mem[4225] = 80'h10100000010000010010;
mem[4226] = 80'h00109400000208004500;
mem[4227] = 80'h0010002e2a740000fffd;
mem[4228] = 80'h00100f06c0550102c000;
mem[4229] = 80'h00100001ffabffabffab;
mem[4230] = 80'h00108b361f70af17d0bb;
mem[4231] = 80'h00106057001589e2efe9;
mem[4232] = 80'h01106e0d8d3f629edcd0;
mem[4233] = 80'h00000000000000000000;
mem[4234] = 80'h00000000000000000000;
mem[4235] = 80'h00000000000000000000;
mem[4236] = 80'h00000000000000000000;
mem[4237] = 80'h10100000010000010010;
mem[4238] = 80'h00109400000208004500;
mem[4239] = 80'h0010002e2a750000fffd;
mem[4240] = 80'h00100f05c0550102c000;
mem[4241] = 80'h00100001ffabffabffab;
mem[4242] = 80'h00108a47c15c776e1204;
mem[4243] = 80'h0010ab8587f87c316fb8;
mem[4244] = 80'h01105d0fae71a42ecf94;
mem[4245] = 80'h00000000000000000000;
mem[4246] = 80'h00000000000000000000;
mem[4247] = 80'h00000000000000000000;
mem[4248] = 80'h10100000010000010010;
mem[4249] = 80'h00109400000208004500;
mem[4250] = 80'h0010002e2a760000fffd;
mem[4251] = 80'h00100f04c0550102c000;
mem[4252] = 80'h00100001ffabffabffab;
mem[4253] = 80'h001089d5a3291fe455c4;
mem[4254] = 80'h0010f7f20fce6241ff4a;
mem[4255] = 80'h0110c79b2c6f31411df5;
mem[4256] = 80'h00000000000000000000;
mem[4257] = 80'h10100000010000010010;
mem[4258] = 80'h00109400000208004500;
mem[4259] = 80'h0010002e2a770000fffd;
mem[4260] = 80'h00100f03c0550102c000;
mem[4261] = 80'h00100001ffabffabffab;
mem[4262] = 80'h001088a47d05c79d977b;
mem[4263] = 80'h00103c2088239791f01b;
mem[4264] = 80'h0110a66fa8dba2e7f98b;
mem[4265] = 80'h00000000000000000000;
mem[4266] = 80'h00000000000000000000;
mem[4267] = 80'h00000000000000000000;
mem[4268] = 80'h00000000000000000000;
mem[4269] = 80'h10100000010000010010;
mem[4270] = 80'h00109400000208004500;
mem[4271] = 80'h0010002e2a780000fffd;
mem[4272] = 80'h00100f02c0550102c000;
mem[4273] = 80'h00100001ffabffabffab;
mem[4274] = 80'h0010879c2afcbdcd4ac5;
mem[4275] = 80'h0010862c2d161b830981;
mem[4276] = 80'h0110d752953abb49985d;
mem[4277] = 80'h00000000000000000000;
mem[4278] = 80'h10100000010000010010;
mem[4279] = 80'h00109400000208004500;
mem[4280] = 80'h0010002e2a790000fffd;
mem[4281] = 80'h00100f01c0550102c000;
mem[4282] = 80'h00100001ffabffabffab;
mem[4283] = 80'h001086edf4d065b4887a;
mem[4284] = 80'h00104dfeaafbee5377d0;
mem[4285] = 80'h01108dcea92506d96e67;
mem[4286] = 80'h00000000000000000000;
mem[4287] = 80'h00000000000000000000;
mem[4288] = 80'h00000000000000000000;
mem[4289] = 80'h00000000000000000000;
mem[4290] = 80'h10100000010000010010;
mem[4291] = 80'h00109400000208004500;
mem[4292] = 80'h0010002e2a7a0000fffd;
mem[4293] = 80'h00100f00c0550102c000;
mem[4294] = 80'h00100001ffabffabffab;
mem[4295] = 80'h0010857f96a50d3ecfba;
mem[4296] = 80'h0010118922cdf0233e22;
mem[4297] = 80'h0110b8e5eb5f0539a269;
mem[4298] = 80'h00000000000000000000;
mem[4299] = 80'h00000000000000000000;
mem[4300] = 80'h00000000000000000000;
mem[4301] = 80'h10100000010000010010;
mem[4302] = 80'h00109400000208004500;
mem[4303] = 80'h0010002e2a7b0000fffd;
mem[4304] = 80'h00100effc0550102c000;
mem[4305] = 80'h00100001ffabffabffab;
mem[4306] = 80'h0010840e4889d5470d05;
mem[4307] = 80'h0010da5ba52005f37773;
mem[4308] = 80'h01107e7bd5bc731d7cc9;
mem[4309] = 80'h00000000000000000000;
mem[4310] = 80'h10100000010000010010;
mem[4311] = 80'h00109400000208004500;
mem[4312] = 80'h0010002e2a7c0000fffd;
mem[4313] = 80'h00100efec0550102c000;
mem[4314] = 80'h00100001ffabffabffab;
mem[4315] = 80'h0010832a8c6304538285;
mem[4316] = 80'h001062b4b44c39125296;
mem[4317] = 80'h0110c23704b86b7e757d;
mem[4318] = 80'h00000000000000000000;
mem[4319] = 80'h00000000000000000000;
mem[4320] = 80'h00000000000000000000;
mem[4321] = 80'h10100000010000010010;
mem[4322] = 80'h00109400000208004500;
mem[4323] = 80'h0010002e2a7d0000fffd;
mem[4324] = 80'h00100efdc0550102c000;
mem[4325] = 80'h00100001ffabffabffab;
mem[4326] = 80'h0010825b524fdc2a403a;
mem[4327] = 80'h0010a96633a1ccc213c7;
mem[4328] = 80'h01108d00c45d31fb24e5;
mem[4329] = 80'h00000000000000000000;
mem[4330] = 80'h00000000000000000000;
mem[4331] = 80'h00000000000000000000;
mem[4332] = 80'h10100000010000010010;
mem[4333] = 80'h00109400000208004500;
mem[4334] = 80'h0010002e2a7e0000fffd;
mem[4335] = 80'h00100efcc0550102c000;
mem[4336] = 80'h00100001ffabffabffab;
mem[4337] = 80'h001081c9303ab4a007fa;
mem[4338] = 80'h0010f511bb97d2b35235;
mem[4339] = 80'h011006b2b51c29a4c3eb;
mem[4340] = 80'h00000000000000000000;
mem[4341] = 80'h10100000010000010010;
mem[4342] = 80'h00109400000208004500;
mem[4343] = 80'h0010002e2a7f0000fffd;
mem[4344] = 80'h00100efbc0550102c000;
mem[4345] = 80'h00100001ffabffabffab;
mem[4346] = 80'h001080b8ee166cd9c545;
mem[4347] = 80'h00103ec33c7a27631264;
mem[4348] = 80'h01107ab42f583c5fe616;
mem[4349] = 80'h00000000000000000000;
mem[4350] = 80'h00000000000000000000;
mem[4351] = 80'h00000000000000000000;
mem[4352] = 80'h00000000000000000000;
mem[4353] = 80'h10100000010000010010;
mem[4354] = 80'h00109400000208004500;
mem[4355] = 80'h0010002e2a800000fffd;
mem[4356] = 80'h00100efac0550102c000;
mem[4357] = 80'h00100001ffabffabffab;
mem[4358] = 80'h00107f97a40ddb0e84d0;
mem[4359] = 80'h001078724121742cd5ab;
mem[4360] = 80'h0110be4fbabf1eb99543;
mem[4361] = 80'h00000000000000000000;
mem[4362] = 80'h00000000000000000000;
mem[4363] = 80'h00000000000000000000;
mem[4364] = 80'h10100000010000010010;
mem[4365] = 80'h00109400000208004500;
mem[4366] = 80'h0010002e2a810000fffd;
mem[4367] = 80'h00100ef9c0550102c000;
mem[4368] = 80'h00100001ffabffabffab;
mem[4369] = 80'h00107ee67a210377466f;
mem[4370] = 80'h0010b3a0c6cc81fcddfa;
mem[4371] = 80'h0110462c9c800ff8a176;
mem[4372] = 80'h00000000000000000000;
mem[4373] = 80'h10100000010000010010;
mem[4374] = 80'h00109400000208004500;
mem[4375] = 80'h0010002e2a820000fffd;
mem[4376] = 80'h00100ef8c0550102c000;
mem[4377] = 80'h00100001ffabffabffab;
mem[4378] = 80'h00107d7418546bfd01af;
mem[4379] = 80'h0010efd74efa9f8c5408;
mem[4380] = 80'h0110655364d07307d3b2;
mem[4381] = 80'h00000000000000000000;
mem[4382] = 80'h00000000000000000000;
mem[4383] = 80'h00000000000000000000;
mem[4384] = 80'h00000000000000000000;
mem[4385] = 80'h10100000010000010010;
mem[4386] = 80'h00109400000208004500;
mem[4387] = 80'h0010002e2a830000fffd;
mem[4388] = 80'h00100ef7c0550102c000;
mem[4389] = 80'h00100001ffabffabffab;
mem[4390] = 80'h00107c05c678b384c310;
mem[4391] = 80'h00102405c9176a5ccd59;
mem[4392] = 80'h0110b6ea6b2e37840a4c;
mem[4393] = 80'h00000000000000000000;
mem[4394] = 80'h00000000000000000000;
mem[4395] = 80'h00000000000000000000;
mem[4396] = 80'h10100000010000010010;
mem[4397] = 80'h00109400000208004500;
mem[4398] = 80'h0010002e2a840000fffd;
mem[4399] = 80'h00100ef6c0550102c000;
mem[4400] = 80'h00100001ffabffabffab;
mem[4401] = 80'h00107b21029262904c90;
mem[4402] = 80'h00109cead87b56bdb6bc;
mem[4403] = 80'h01102716293577d3e58e;
mem[4404] = 80'h00000000000000000000;
mem[4405] = 80'h00000000000000000000;
mem[4406] = 80'h00000000000000000000;
mem[4407] = 80'h10100000010000010010;
mem[4408] = 80'h00109400000208004500;
mem[4409] = 80'h0010002e2a850000fffd;
mem[4410] = 80'h00100ef5c0550102c000;
mem[4411] = 80'h00100001ffabffabffab;
mem[4412] = 80'h00107a50dcbebae98e2f;
mem[4413] = 80'h001057385f96a36db9ed;
mem[4414] = 80'h011046e204cb68895791;
mem[4415] = 80'h00000000000000000000;
mem[4416] = 80'h10100000010000010010;
mem[4417] = 80'h00109400000208004500;
mem[4418] = 80'h0010002e2a860000fffd;
mem[4419] = 80'h00100ef4c0550102c000;
mem[4420] = 80'h00100001ffabffabffab;
mem[4421] = 80'h001079c2becbd263c9ef;
mem[4422] = 80'h00100b4fd7a0bd1d0a1f;
mem[4423] = 80'h01108fc3f12dcd9888b8;
mem[4424] = 80'h00000000000000000000;
mem[4425] = 80'h00000000000000000000;
mem[4426] = 80'h00000000000000000000;
mem[4427] = 80'h10100000010000010010;
mem[4428] = 80'h00109400000208004500;
mem[4429] = 80'h0010002e2a870000fffd;
mem[4430] = 80'h00100ef3c0550102c000;
mem[4431] = 80'h00100001ffabffabffab;
mem[4432] = 80'h001078b360e70a1a0b50;
mem[4433] = 80'h0010c09d504d48cd494e;
mem[4434] = 80'h0110a696c75d5f791672;
mem[4435] = 80'h00000000000000000000;
mem[4436] = 80'h00000000000000000000;
mem[4437] = 80'h00000000000000000000;
mem[4438] = 80'h10100000010000010010;
mem[4439] = 80'h00109400000208004500;
mem[4440] = 80'h0010002e2a880000fffd;
mem[4441] = 80'h00100ef2c0550102c000;
mem[4442] = 80'h00100001ffabffabffab;
mem[4443] = 80'h0010778b371e704ad6ee;
mem[4444] = 80'h00107a91f578c4d87fd4;
mem[4445] = 80'h011054510114d6b994e9;
mem[4446] = 80'h00000000000000000000;
mem[4447] = 80'h00000000000000000000;
mem[4448] = 80'h00000000000000000000;
mem[4449] = 80'h10100000010000010010;
mem[4450] = 80'h00109400000208004500;
mem[4451] = 80'h0010002e2a890000fffd;
mem[4452] = 80'h00100ef1c0550102c000;
mem[4453] = 80'h00100001ffabffabffab;
mem[4454] = 80'h001076fae932a8331451;
mem[4455] = 80'h0010b143729531082085;
mem[4456] = 80'h01103b1a32cd94af3ea5;
mem[4457] = 80'h00000000000000000000;
mem[4458] = 80'h10100000010000010010;
mem[4459] = 80'h00109400000208004500;
mem[4460] = 80'h0010002e2a8a0000fffd;
mem[4461] = 80'h00100ef0c0550102c000;
mem[4462] = 80'h00100001ffabffabffab;
mem[4463] = 80'h001075688b47c0b95391;
mem[4464] = 80'h0010ed34faa32f78e877;
mem[4465] = 80'h01102698c4a315d64257;
mem[4466] = 80'h00000000000000000000;
mem[4467] = 80'h00000000000000000000;
mem[4468] = 80'h00000000000000000000;
mem[4469] = 80'h10100000010000010010;
mem[4470] = 80'h00109400000208004500;
mem[4471] = 80'h0010002e2a8b0000fffd;
mem[4472] = 80'h00100eefc0550102c000;
mem[4473] = 80'h00100001ffabffabffab;
mem[4474] = 80'h00107419556b18c0912e;
mem[4475] = 80'h001026e67d4edaa8a026;
mem[4476] = 80'h0110d3379a5018e1e07f;
mem[4477] = 80'h00000000000000000000;
mem[4478] = 80'h00000000000000000000;
mem[4479] = 80'h00000000000000000000;
mem[4480] = 80'h10100000010000010010;
mem[4481] = 80'h00109400000208004500;
mem[4482] = 80'h0010002e2a8c0000fffd;
mem[4483] = 80'h00100eeec0550102c000;
mem[4484] = 80'h00100001ffabffabffab;
mem[4485] = 80'h0010733d9181c9d41eae;
mem[4486] = 80'h00109e096c22e649e4c3;
mem[4487] = 80'h01105760e6231be465f8;
mem[4488] = 80'h00000000000000000000;
mem[4489] = 80'h00000000000000000000;
mem[4490] = 80'h00000000000000000000;
mem[4491] = 80'h10100000010000010010;
mem[4492] = 80'h00109400000208004500;
mem[4493] = 80'h0010002e2a8d0000fffd;
mem[4494] = 80'h00100eedc0550102c000;
mem[4495] = 80'h00100001ffabffabffab;
mem[4496] = 80'h0010724c4fad11addc11;
mem[4497] = 80'h001055dbebcf13996792;
mem[4498] = 80'h011068612b0f19e3db20;
mem[4499] = 80'h00000000000000000000;
mem[4500] = 80'h10100000010000010010;
mem[4501] = 80'h00109400000208004500;
mem[4502] = 80'h0010002e2a8e0000fffd;
mem[4503] = 80'h00100eecc0550102c000;
mem[4504] = 80'h00100001ffabffabffab;
mem[4505] = 80'h001071de2dd879279bd1;
mem[4506] = 80'h001009ac63f90de9e460;
mem[4507] = 80'h0110a4d5468b5e7f5cdb;
mem[4508] = 80'h00000000000000000000;
mem[4509] = 80'h00000000000000000000;
mem[4510] = 80'h00000000000000000000;
mem[4511] = 80'h10100000010000010010;
mem[4512] = 80'h00109400000208004500;
mem[4513] = 80'h0010002e2a8f0000fffd;
mem[4514] = 80'h00100eebc0550102c000;
mem[4515] = 80'h00100001ffabffabffab;
mem[4516] = 80'h001070aff3f4a15e596e;
mem[4517] = 80'h0010c27ee414f839fb31;
mem[4518] = 80'h0110c652403cc209d072;
mem[4519] = 80'h00000000000000000000;
mem[4520] = 80'h00000000000000000000;
mem[4521] = 80'h00000000000000000000;
mem[4522] = 80'h00000000000000000000;
mem[4523] = 80'h10100000010000010010;
mem[4524] = 80'h00109400000208004500;
mem[4525] = 80'h0010002e2a900000fffd;
mem[4526] = 80'h00100eeac0550102c000;
mem[4527] = 80'h00100001ffabffabffab;
mem[4528] = 80'h00106fae822a8d8620ac;
mem[4529] = 80'h00107db5299215cc0f54;
mem[4530] = 80'h0110cc75c71623a87c75;
mem[4531] = 80'h00000000000000000000;
mem[4532] = 80'h10100000010000010010;
mem[4533] = 80'h00109400000208004500;
mem[4534] = 80'h0010002e2a910000fffd;
mem[4535] = 80'h00100ee9c0550102c000;
mem[4536] = 80'h00100001ffabffabffab;
mem[4537] = 80'h00106edf5c0655ffe213;
mem[4538] = 80'h0010b667ae7fe01d8605;
mem[4539] = 80'h01102b8f066def01e5a9;
mem[4540] = 80'h00000000000000000000;
mem[4541] = 80'h00000000000000000000;
mem[4542] = 80'h00000000000000000000;
mem[4543] = 80'h10100000010000010010;
mem[4544] = 80'h00109400000208004500;
mem[4545] = 80'h0010002e2a920000fffd;
mem[4546] = 80'h00100ee8c0550102c000;
mem[4547] = 80'h00100001ffabffabffab;
mem[4548] = 80'h00106d4d3e733d75a5d3;
mem[4549] = 80'h0010ea102649fe6d0ff7;
mem[4550] = 80'h011008f04947ce5ec376;
mem[4551] = 80'h00000000000000000000;
mem[4552] = 80'h00000000000000000000;
mem[4553] = 80'h00000000000000000000;
mem[4554] = 80'h10100000010000010010;
mem[4555] = 80'h00109400000208004500;
mem[4556] = 80'h0010002e2a930000fffd;
mem[4557] = 80'h00100ee7c0550102c000;
mem[4558] = 80'h00100001ffabffabffab;
mem[4559] = 80'h00106c3ce05fe50c676c;
mem[4560] = 80'h001021c2a1a40bbd77a6;
mem[4561] = 80'h0110f8ca27551144acd1;
mem[4562] = 80'h00000000000000000000;
mem[4563] = 80'h00000000000000000000;
mem[4564] = 80'h00000000000000000000;
mem[4565] = 80'h10100000010000010010;
mem[4566] = 80'h00109400000208004500;
mem[4567] = 80'h0010002e2a940000fffd;
mem[4568] = 80'h00100ee6c0550102c000;
mem[4569] = 80'h00100001ffabffabffab;
mem[4570] = 80'h00106b1824b53418e8ec;
mem[4571] = 80'h0010992db0c8375c4343;
mem[4572] = 80'h011074c419d3175a4af4;
mem[4573] = 80'h00000000000000000000;
mem[4574] = 80'h10100000010000010010;
mem[4575] = 80'h00109400000208004500;
mem[4576] = 80'h0010002e2a950000fffd;
mem[4577] = 80'h00100ee5c0550102c000;
mem[4578] = 80'h00100001ffabffabffab;
mem[4579] = 80'h00106a69fa99ec612a53;
mem[4580] = 80'h001052ff3725c28c0312;
mem[4581] = 80'h011008c22bc23a612afc;
mem[4582] = 80'h00000000000000000000;
mem[4583] = 80'h00000000000000000000;
mem[4584] = 80'h00000000000000000000;
mem[4585] = 80'h10100000010000010010;
mem[4586] = 80'h00109400000208004500;
mem[4587] = 80'h0010002e2a960000fffd;
mem[4588] = 80'h00100ee4c0550102c000;
mem[4589] = 80'h00100001ffabffabffab;
mem[4590] = 80'h001069fb98ec84eb6d93;
mem[4591] = 80'h00100e88bf13dcfc52e0;
mem[4592] = 80'h0110b73355ec640b6c00;
mem[4593] = 80'h00000000000000000000;
mem[4594] = 80'h00000000000000000000;
mem[4595] = 80'h00000000000000000000;
mem[4596] = 80'h10100000010000010010;
mem[4597] = 80'h00109400000208004500;
mem[4598] = 80'h0010002e2a970000fffd;
mem[4599] = 80'h00100ee3c0550102c000;
mem[4600] = 80'h00100001ffabffabffab;
mem[4601] = 80'h0010688a46c05c92af2c;
mem[4602] = 80'h0010c55a38fe292c13b1;
mem[4603] = 80'h0110f80411bb7352276a;
mem[4604] = 80'h00000000000000000000;
mem[4605] = 80'h00000000000000000000;
mem[4606] = 80'h00000000000000000000;
mem[4607] = 80'h10100000010000010010;
mem[4608] = 80'h00109400000208004500;
mem[4609] = 80'h0010002e2a980000fffd;
mem[4610] = 80'h00100ee2c0550102c000;
mem[4611] = 80'h00100001ffabffabffab;
mem[4612] = 80'h001067b2113926c27292;
mem[4613] = 80'h00107f569dcba53ea32b;
mem[4614] = 80'h01103e6d49c60c17329e;
mem[4615] = 80'h00000000000000000000;
mem[4616] = 80'h10100000010000010010;
mem[4617] = 80'h00109400000208004500;
mem[4618] = 80'h0010002e2a990000fffd;
mem[4619] = 80'h00100ee1c0550102c000;
mem[4620] = 80'h00100001ffabffabffab;
mem[4621] = 80'h001066c3cf15febbb02d;
mem[4622] = 80'h0010b4841a2650eeda7a;
mem[4623] = 80'h0110fd6623c26c8451e7;
mem[4624] = 80'h00000000000000000000;
mem[4625] = 80'h00000000000000000000;
mem[4626] = 80'h00000000000000000000;
mem[4627] = 80'h10100000010000010010;
mem[4628] = 80'h00109400000208004500;
mem[4629] = 80'h0010002e2a9a0000fffd;
mem[4630] = 80'h00100ee0c0550102c000;
mem[4631] = 80'h00100001ffabffabffab;
mem[4632] = 80'h00106551ad609631f7ed;
mem[4633] = 80'h0010e8f392104e9e5388;
mem[4634] = 80'h0110de1963e914f7e8c8;
mem[4635] = 80'h00000000000000000000;
mem[4636] = 80'h00000000000000000000;
mem[4637] = 80'h00000000000000000000;
mem[4638] = 80'h10100000010000010010;
mem[4639] = 80'h00109400000208004500;
mem[4640] = 80'h0010002e2a9b0000fffd;
mem[4641] = 80'h00100edfc0550102c000;
mem[4642] = 80'h00100001ffabffabffab;
mem[4643] = 80'h00106420734c4e483552;
mem[4644] = 80'h0010232115fdbb4ddad9;
mem[4645] = 80'h011057837e2fb97f4c1a;
mem[4646] = 80'h00000000000000000000;
mem[4647] = 80'h00000000000000000000;
mem[4648] = 80'h00000000000000000000;
mem[4649] = 80'h10100000010000010010;
mem[4650] = 80'h00109400000208004500;
mem[4651] = 80'h0010002e2a9c0000fffd;
mem[4652] = 80'h00100edec0550102c000;
mem[4653] = 80'h00100001ffabffabffab;
mem[4654] = 80'h00106304b7a69f5cbad2;
mem[4655] = 80'h00109bce049187aca13c;
mem[4656] = 80'h0110c67ffb5c1a80711f;
mem[4657] = 80'h00000000000000000000;
mem[4658] = 80'h10100000010000010010;
mem[4659] = 80'h00109400000208004500;
mem[4660] = 80'h0010002e2a9d0000fffd;
mem[4661] = 80'h00100eddc0550102c000;
mem[4662] = 80'h00100001ffabffabffab;
mem[4663] = 80'h00106275698a4725786d;
mem[4664] = 80'h0010501c837c727cbe6d;
mem[4665] = 80'h0110a4f8caf16afc0253;
mem[4666] = 80'h00000000000000000000;
mem[4667] = 80'h00000000000000000000;
mem[4668] = 80'h00000000000000000000;
mem[4669] = 80'h00000000000000000000;
mem[4670] = 80'h10100000010000010010;
mem[4671] = 80'h00109400000208004500;
mem[4672] = 80'h0010002e2a9e0000fffd;
mem[4673] = 80'h00100edcc0550102c000;
mem[4674] = 80'h00100001ffabffabffab;
mem[4675] = 80'h001061e70bff2faf3fad;
mem[4676] = 80'h00100c6b0b4a6c0c3e9f;
mem[4677] = 80'h01103d1f233d17e9d09b;
mem[4678] = 80'h00000000000000000000;
mem[4679] = 80'h00000000000000000000;
mem[4680] = 80'h00000000000000000000;
mem[4681] = 80'h10100000010000010010;
mem[4682] = 80'h00109400000208004500;
mem[4683] = 80'h0010002e2a9f0000fffd;
mem[4684] = 80'h00100edbc0550102c000;
mem[4685] = 80'h00100001ffabffabffab;
mem[4686] = 80'h00106096d5d3f7d6fd12;
mem[4687] = 80'h0010c7b98ca799dcbece;
mem[4688] = 80'h0110574dd0518dfa50e8;
mem[4689] = 80'h00000000000000000000;
mem[4690] = 80'h10100000010000010010;
mem[4691] = 80'h00109400000208004500;
mem[4692] = 80'h0010002e2aa00000fffd;
mem[4693] = 80'h00100edac0550102c000;
mem[4694] = 80'h00100001ffabffabffab;
mem[4695] = 80'h00105fe5e843761fcc28;
mem[4696] = 80'h001073fc9047b7e76055;
mem[4697] = 80'h01109dfabb129c428ec4;
mem[4698] = 80'h00000000000000000000;
mem[4699] = 80'h00000000000000000000;
mem[4700] = 80'h00000000000000000000;
mem[4701] = 80'h10100000010000010010;
mem[4702] = 80'h00109400000208004500;
mem[4703] = 80'h0010002e2aa10000fffd;
mem[4704] = 80'h00100ed9c0550102c000;
mem[4705] = 80'h00100001ffabffabffab;
mem[4706] = 80'h00105e94366fae660e97;
mem[4707] = 80'h0010b82e17aa42372b04;
mem[4708] = 80'h01103d0633e4bc48bc52;
mem[4709] = 80'h00000000000000000000;
mem[4710] = 80'h00000000000000000000;
mem[4711] = 80'h00000000000000000000;
mem[4712] = 80'h10100000010000010010;
mem[4713] = 80'h00109400000208004500;
mem[4714] = 80'h0010002e2aa20000fffd;
mem[4715] = 80'h00100ed8c0550102c000;
mem[4716] = 80'h00100001ffabffabffab;
mem[4717] = 80'h00105d06541ac6ec4957;
mem[4718] = 80'h0010e4599f9c5c47e0f6;
mem[4719] = 80'h011075d7078fa96ddb3d;
mem[4720] = 80'h00000000000000000000;
mem[4721] = 80'h00000000000000000000;
mem[4722] = 80'h00000000000000000000;
mem[4723] = 80'h10100000010000010010;
mem[4724] = 80'h00109400000208004500;
mem[4725] = 80'h0010002e2aa30000fffd;
mem[4726] = 80'h00100ed7c0550102c000;
mem[4727] = 80'h00100001ffabffabffab;
mem[4728] = 80'h00105c778a361e958be8;
mem[4729] = 80'h00102f8b1871a997bfa7;
mem[4730] = 80'h01101a9ca2fc26eeb622;
mem[4731] = 80'h00000000000000000000;
mem[4732] = 80'h10100000010000010010;
mem[4733] = 80'h00109400000208004500;
mem[4734] = 80'h0010002e2aa40000fffd;
mem[4735] = 80'h00100ed6c0550102c000;
mem[4736] = 80'h00100001ffabffabffab;
mem[4737] = 80'h00105b534edccf810468;
mem[4738] = 80'h00109764091d95770c42;
mem[4739] = 80'h011023ad1bfe448a1e39;
mem[4740] = 80'h00000000000000000000;
mem[4741] = 80'h00000000000000000000;
mem[4742] = 80'h00000000000000000000;
mem[4743] = 80'h10100000010000010010;
mem[4744] = 80'h00109400000208004500;
mem[4745] = 80'h0010002e2aa50000fffd;
mem[4746] = 80'h00100ed5c0550102c000;
mem[4747] = 80'h00100001ffabffabffab;
mem[4748] = 80'h00105a2290f017f8c6d7;
mem[4749] = 80'h00105cb68ef060a74f13;
mem[4750] = 80'h01100af88fc332db46ef;
mem[4751] = 80'h00000000000000000000;
mem[4752] = 80'h00000000000000000000;
mem[4753] = 80'h00000000000000000000;
mem[4754] = 80'h10100000010000010010;
mem[4755] = 80'h00109400000208004500;
mem[4756] = 80'h0010002e2aa60000fffd;
mem[4757] = 80'h00100ed4c0550102c000;
mem[4758] = 80'h00100001ffabffabffab;
mem[4759] = 80'h001059b0f2857f728117;
mem[4760] = 80'h001000c106c67ed7fde1;
mem[4761] = 80'h0110f0e83e16cd2a37e1;
mem[4762] = 80'h00000000000000000000;
mem[4763] = 80'h00000000000000000000;
mem[4764] = 80'h00000000000000000000;
mem[4765] = 80'h10100000010000010010;
mem[4766] = 80'h00109400000208004500;
mem[4767] = 80'h0010002e2aa70000fffd;
mem[4768] = 80'h00100ed3c0550102c000;
mem[4769] = 80'h00100001ffabffabffab;
mem[4770] = 80'h001058c12ca9a70b43a8;
mem[4771] = 80'h0010cb13812b8b07fdb0;
mem[4772] = 80'h0110812239c7d1ff1f3d;
mem[4773] = 80'h00000000000000000000;
mem[4774] = 80'h10100000010000010010;
mem[4775] = 80'h00109400000208004500;
mem[4776] = 80'h0010002e2aa80000fffd;
mem[4777] = 80'h00100ed2c0550102c000;
mem[4778] = 80'h00100001ffabffabffab;
mem[4779] = 80'h001057f97b50dd5b9e16;
mem[4780] = 80'h0010711f241e07150d2a;
mem[4781] = 80'h01104a87bd3f87fad21c;
mem[4782] = 80'h00000000000000000000;
mem[4783] = 80'h00000000000000000000;
mem[4784] = 80'h00000000000000000000;
mem[4785] = 80'h00000000000000000000;
mem[4786] = 80'h10100000010000010010;
mem[4787] = 80'h00109400000208004500;
mem[4788] = 80'h0010002e2aa90000fffd;
mem[4789] = 80'h00100ed1c0550102c000;
mem[4790] = 80'h00100001ffabffabffab;
mem[4791] = 80'h00105688a57c05225ca9;
mem[4792] = 80'h0010bacda3f3f2c5957b;
mem[4793] = 80'h0110aa0f111dfcf1f0a6;
mem[4794] = 80'h00000000000000000000;
mem[4795] = 80'h00000000000000000000;
mem[4796] = 80'h00000000000000000000;
mem[4797] = 80'h10100000010000010010;
mem[4798] = 80'h00109400000208004500;
mem[4799] = 80'h0010002e2aaa0000fffd;
mem[4800] = 80'h00100ed0c0550102c000;
mem[4801] = 80'h00100001ffabffabffab;
mem[4802] = 80'h0010551ac7096da81b69;
mem[4803] = 80'h0010e6ba2bc5ecb51d89;
mem[4804] = 80'h0110ba4183c9d9c12e1b;
mem[4805] = 80'h00000000000000000000;
mem[4806] = 80'h10100000010000010010;
mem[4807] = 80'h00109400000208004500;
mem[4808] = 80'h0010002e2aab0000fffd;
mem[4809] = 80'h00100ecfc0550102c000;
mem[4810] = 80'h00100001ffabffabffab;
mem[4811] = 80'h0010546b1925b5d1d9d6;
mem[4812] = 80'h00102d68ac28196515d8;
mem[4813] = 80'h01104222b7d63f66a560;
mem[4814] = 80'h00000000000000000000;
mem[4815] = 80'h00000000000000000000;
mem[4816] = 80'h00000000000000000000;
mem[4817] = 80'h10100000010000010010;
mem[4818] = 80'h00109400000208004500;
mem[4819] = 80'h0010002e2aac0000fffd;
mem[4820] = 80'h00100ecec0550102c000;
mem[4821] = 80'h00100001ffabffabffab;
mem[4822] = 80'h0010534fddcf64c55656;
mem[4823] = 80'h00109587bd442584503d;
mem[4824] = 80'h0110f54455f2b20b86f1;
mem[4825] = 80'h00000000000000000000;
mem[4826] = 80'h00000000000000000000;
mem[4827] = 80'h00000000000000000000;
mem[4828] = 80'h10100000010000010010;
mem[4829] = 80'h00109400000208004500;
mem[4830] = 80'h0010002e2aad0000fffd;
mem[4831] = 80'h00100ecdc0550102c000;
mem[4832] = 80'h00100001ffabffabffab;
mem[4833] = 80'h0010523e03e3bcbc94e9;
mem[4834] = 80'h00105e553aa9d054116c;
mem[4835] = 80'h0110ba7323059ef6f128;
mem[4836] = 80'h00000000000000000000;
mem[4837] = 80'h00000000000000000000;
mem[4838] = 80'h00000000000000000000;
mem[4839] = 80'h10100000010000010010;
mem[4840] = 80'h00109400000208004500;
mem[4841] = 80'h0010002e2aae0000fffd;
mem[4842] = 80'h00100eccc0550102c000;
mem[4843] = 80'h00100001ffabffabffab;
mem[4844] = 80'h001051ac6196d436d329;
mem[4845] = 80'h00100222b29fce3b509e;
mem[4846] = 80'h011069a3681d3f410363;
mem[4847] = 80'h00000000000000000000;
mem[4848] = 80'h10100000010000010010;
mem[4849] = 80'h00109400000208004500;
mem[4850] = 80'h0010002e2aaf0000fffd;
mem[4851] = 80'h00100ecbc0550102c000;
mem[4852] = 80'h00100001ffabffabffab;
mem[4853] = 80'h001050ddbfba0c4f1196;
mem[4854] = 80'h0010c9f035723beb11cf;
mem[4855] = 80'h011026945dd1531ab158;
mem[4856] = 80'h00000000000000000000;
mem[4857] = 80'h00000000000000000000;
mem[4858] = 80'h00000000000000000000;
mem[4859] = 80'h10100000010000010010;
mem[4860] = 80'h00109400000208004500;
mem[4861] = 80'h0010002e2ab00000fffd;
mem[4862] = 80'h00100ecac0550102c000;
mem[4863] = 80'h00100001ffabffabffab;
mem[4864] = 80'h00104fdcce6420976854;
mem[4865] = 80'h0010763bf8f4d61ebbaa;
mem[4866] = 80'h0110010356d6f4d0762c;
mem[4867] = 80'h00000000000000000000;
mem[4868] = 80'h00000000000000000000;
mem[4869] = 80'h00000000000000000000;
mem[4870] = 80'h10100000010000010010;
mem[4871] = 80'h00109400000208004500;
mem[4872] = 80'h0010002e2ab10000fffd;
mem[4873] = 80'h00100ec9c0550102c000;
mem[4874] = 80'h00100001ffabffabffab;
mem[4875] = 80'h00104ead1048f8eeaaeb;
mem[4876] = 80'h0010bde97f1923cef1fb;
mem[4877] = 80'h011092ce17940bca1b60;
mem[4878] = 80'h00000000000000000000;
mem[4879] = 80'h00000000000000000000;
mem[4880] = 80'h00000000000000000000;
mem[4881] = 80'h10100000010000010010;
mem[4882] = 80'h00109400000208004500;
mem[4883] = 80'h0010002e2ab20000fffd;
mem[4884] = 80'h00100ec8c0550102c000;
mem[4885] = 80'h00100001ffabffabffab;
mem[4886] = 80'h00104d3f723d9064ed2b;
mem[4887] = 80'h0010e19ef72f3dbebb09;
mem[4888] = 80'h0110f2b6fea473fa90a1;
mem[4889] = 80'h00000000000000000000;
mem[4890] = 80'h10100000010000010010;
mem[4891] = 80'h00109400000208004500;
mem[4892] = 80'h0010002e2ab30000fffd;
mem[4893] = 80'h00100ec7c0550102c000;
mem[4894] = 80'h00100001ffabffabffab;
mem[4895] = 80'h00104c4eac11481d2f94;
mem[4896] = 80'h00102a4c70c2c86ec258;
mem[4897] = 80'h011031bd385bc543f1b2;
mem[4898] = 80'h00000000000000000000;
mem[4899] = 80'h00000000000000000000;
mem[4900] = 80'h00000000000000000000;
mem[4901] = 80'h00000000000000000000;
mem[4902] = 80'h10100000010000010010;
mem[4903] = 80'h00109400000208004500;
mem[4904] = 80'h0010002e2ab40000fffd;
mem[4905] = 80'h00100ec6c0550102c000;
mem[4906] = 80'h00100001ffabffabffab;
mem[4907] = 80'h00104b6a68fb9909a014;
mem[4908] = 80'h001092a361aef48fb6bd;
mem[4909] = 80'h0110b07fc25caa41b9c7;
mem[4910] = 80'h00000000000000000000;
mem[4911] = 80'h00000000000000000000;
mem[4912] = 80'h00000000000000000000;
mem[4913] = 80'h10100000010000010010;
mem[4914] = 80'h00109400000208004500;
mem[4915] = 80'h0010002e2ab50000fffd;
mem[4916] = 80'h00100ec5c0550102c000;
mem[4917] = 80'h00100001ffabffabffab;
mem[4918] = 80'h00104a1bb6d7417062ab;
mem[4919] = 80'h00105971e643015fb6ec;
mem[4920] = 80'h0110c1b5a13a984f9fc7;
mem[4921] = 80'h00000000000000000000;
mem[4922] = 80'h10100000010000010010;
mem[4923] = 80'h00109400000208004500;
mem[4924] = 80'h0010002e2ab60000fffd;
mem[4925] = 80'h00100ec4c0550102c000;
mem[4926] = 80'h00100001ffabffabffab;
mem[4927] = 80'h00104989d4a229fa256b;
mem[4928] = 80'h001005066e751f2f261e;
mem[4929] = 80'h01105b217e84fca08e7f;
mem[4930] = 80'h00000000000000000000;
mem[4931] = 80'h00000000000000000000;
mem[4932] = 80'h00000000000000000000;
mem[4933] = 80'h10100000010000010010;
mem[4934] = 80'h00109400000208004500;
mem[4935] = 80'h0010002e2ab70000fffd;
mem[4936] = 80'h00100ec3c0550102c000;
mem[4937] = 80'h00100001ffabffabffab;
mem[4938] = 80'h001048f80a8ef183e7d4;
mem[4939] = 80'h0010ced4e998eafea94f;
mem[4940] = 80'h0110167d6fe7753ca390;
mem[4941] = 80'h00000000000000000000;
mem[4942] = 80'h00000000000000000000;
mem[4943] = 80'h00000000000000000000;
mem[4944] = 80'h10100000010000010010;
mem[4945] = 80'h00109400000208004500;
mem[4946] = 80'h0010002e2ab80000fffd;
mem[4947] = 80'h00100ec2c0550102c000;
mem[4948] = 80'h00100001ffabffabffab;
mem[4949] = 80'h001047c05d778bd33a6a;
mem[4950] = 80'h001074d84cad66ec57d5;
mem[4951] = 80'h0110fed7156ba866e8ef;
mem[4952] = 80'h00000000000000000000;
mem[4953] = 80'h00000000000000000000;
mem[4954] = 80'h00000000000000000000;
mem[4955] = 80'h10100000010000010010;
mem[4956] = 80'h00109400000208004500;
mem[4957] = 80'h0010002e2ab90000fffd;
mem[4958] = 80'h00100ec1c0550102c000;
mem[4959] = 80'h00100001ffabffabffab;
mem[4960] = 80'h001046b1835b53aaf8d5;
mem[4961] = 80'h0010bf0acb40933c2c84;
mem[4962] = 80'h01105bbe43a8becdaef8;
mem[4963] = 80'h00000000000000000000;
mem[4964] = 80'h10100000010000010010;
mem[4965] = 80'h00109400000208004500;
mem[4966] = 80'h0010002e2aba0000fffd;
mem[4967] = 80'h00100ec0c0550102c000;
mem[4968] = 80'h00100001ffabffabffab;
mem[4969] = 80'h00104523e12e3b20bf15;
mem[4970] = 80'h0010e37d43768d4ce776;
mem[4971] = 80'h0110136f305101c3f036;
mem[4972] = 80'h00000000000000000000;
mem[4973] = 80'h00000000000000000000;
mem[4974] = 80'h00000000000000000000;
mem[4975] = 80'h10100000010000010010;
mem[4976] = 80'h00109400000208004500;
mem[4977] = 80'h0010002e2abb0000fffd;
mem[4978] = 80'h00100ebfc0550102c000;
mem[4979] = 80'h00100001ffabffabffab;
mem[4980] = 80'h001044523f02e3597daa;
mem[4981] = 80'h001028afc49b789ca827;
mem[4982] = 80'h01107f578e40ac2b5550;
mem[4983] = 80'h00000000000000000000;
mem[4984] = 80'h00000000000000000000;
mem[4985] = 80'h00000000000000000000;
mem[4986] = 80'h10100000010000010010;
mem[4987] = 80'h00109400000208004500;
mem[4988] = 80'h0010002e2abc0000fffd;
mem[4989] = 80'h00100ebec0550102c000;
mem[4990] = 80'h00100001ffabffabffab;
mem[4991] = 80'h00104376fbe8324df22a;
mem[4992] = 80'h00109040d5f7447d0ac2;
mem[4993] = 80'h01104114a59c8806becd;
mem[4994] = 80'h00000000000000000000;
mem[4995] = 80'h00000000000000000000;
mem[4996] = 80'h00000000000000000000;
mem[4997] = 80'h10100000010000010010;
mem[4998] = 80'h00109400000208004500;
mem[4999] = 80'h0010002e2abd0000fffd;
mem[5000] = 80'h00100ebdc0550102c000;
mem[5001] = 80'h00100001ffabffabffab;
mem[5002] = 80'h0010420725c4ea343095;
mem[5003] = 80'h00105b92521ab1ad4893;
mem[5004] = 80'h01105b707a0c281567ac;
mem[5005] = 80'h00000000000000000000;
mem[5006] = 80'h10100000010000010010;
mem[5007] = 80'h00109400000208004500;
mem[5008] = 80'h0010002e2abe0000fffd;
mem[5009] = 80'h00100ebcc0550102c000;
mem[5010] = 80'h00100001ffabffabffab;
mem[5011] = 80'h0010419547b182be7755;
mem[5012] = 80'h001007e5da2cafdd8a61;
mem[5013] = 80'h0110a939b71a36710a8e;
mem[5014] = 80'h00000000000000000000;
mem[5015] = 80'h00000000000000000000;
mem[5016] = 80'h00000000000000000000;
mem[5017] = 80'h10100000010000010010;
mem[5018] = 80'h00109400000208004500;
mem[5019] = 80'h0010002e2abf0000fffd;
mem[5020] = 80'h00100ebbc0550102c000;
mem[5021] = 80'h00100001ffabffabffab;
mem[5022] = 80'h001040e4999d5ac7b5ea;
mem[5023] = 80'h0010cc375dc15a0dcb30;
mem[5024] = 80'h0110e60edf850d09cf48;
mem[5025] = 80'h00000000000000000000;
mem[5026] = 80'h00000000000000000000;
mem[5027] = 80'h00000000000000000000;
mem[5028] = 80'h10100000010000010010;
mem[5029] = 80'h00109400000208004500;
mem[5030] = 80'h0010002e2ac00000fffd;
mem[5031] = 80'h00100ebac0550102c000;
mem[5032] = 80'h00100001ffabffabffab;
mem[5033] = 80'h00103f733c90812c1520;
mem[5034] = 80'h00106f6fe3ecf3aa3e57;
mem[5035] = 80'h011096eed1622dce5915;
mem[5036] = 80'h00000000000000000000;
mem[5037] = 80'h00000000000000000000;
mem[5038] = 80'h00000000000000000000;
mem[5039] = 80'h10100000010000010010;
mem[5040] = 80'h00109400000208004500;
mem[5041] = 80'h0010002e2ac10000fffd;
mem[5042] = 80'h00100eb9c0550102c000;
mem[5043] = 80'h00100001ffabffabffab;
mem[5044] = 80'h00103e02e2bc5955d79f;
mem[5045] = 80'h0010a4bd64010679b606;
mem[5046] = 80'h01102c45bcc7a33ac3a2;
mem[5047] = 80'h00000000000000000000;
mem[5048] = 80'h10100000010000010010;
mem[5049] = 80'h00109400000208004500;
mem[5050] = 80'h0010002e2ac20000fffd;
mem[5051] = 80'h00100eb8c0550102c000;
mem[5052] = 80'h00100001ffabffabffab;
mem[5053] = 80'h00103d9080c931df905f;
mem[5054] = 80'h0010f8caec3718093ff4;
mem[5055] = 80'h01100f3a332d7c707b2d;
mem[5056] = 80'h00000000000000000000;
mem[5057] = 80'h00000000000000000000;
mem[5058] = 80'h00000000000000000000;
mem[5059] = 80'h00000000000000000000;
mem[5060] = 80'h10100000010000010010;
mem[5061] = 80'h00109400000208004500;
mem[5062] = 80'h0010002e2ac30000fffd;
mem[5063] = 80'h00100eb7c0550102c000;
mem[5064] = 80'h00100001ffabffabffab;
mem[5065] = 80'h00103ce15ee5e9a652e0;
mem[5066] = 80'h001033186bdaedd926a5;
mem[5067] = 80'h0110c71bad24d20289f2;
mem[5068] = 80'h00000000000000000000;
mem[5069] = 80'h00000000000000000000;
mem[5070] = 80'h00000000000000000000;
mem[5071] = 80'h10100000010000010010;
mem[5072] = 80'h00109400000208004500;
mem[5073] = 80'h0010002e2ac40000fffd;
mem[5074] = 80'h00100eb6c0550102c000;
mem[5075] = 80'h00100001ffabffabffab;
mem[5076] = 80'h00103bc59a0f38b2dd60;
mem[5077] = 80'h00108bf77ab6d1385340;
mem[5078] = 80'h011075e873081613fed6;
mem[5079] = 80'h00000000000000000000;
mem[5080] = 80'h10100000010000010010;
mem[5081] = 80'h00109400000208004500;
mem[5082] = 80'h0010002e2ac50000fffd;
mem[5083] = 80'h00100eb5c0550102c000;
mem[5084] = 80'h00100001ffabffabffab;
mem[5085] = 80'h00103ab44423e0cb1fdf;
mem[5086] = 80'h00104025fd5b24e8d211;
mem[5087] = 80'h01102c8b1f77688fe853;
mem[5088] = 80'h00000000000000000000;
mem[5089] = 80'h00000000000000000000;
mem[5090] = 80'h00000000000000000000;
mem[5091] = 80'h10100000010000010010;
mem[5092] = 80'h00109400000208004500;
mem[5093] = 80'h0010002e2ac60000fffd;
mem[5094] = 80'h00100eb4c0550102c000;
mem[5095] = 80'h00100001ffabffabffab;
mem[5096] = 80'h0010392626568841581f;
mem[5097] = 80'h00101c52756d3a9863e3;
mem[5098] = 80'h011083c80c1f1a72c560;
mem[5099] = 80'h00000000000000000000;
mem[5100] = 80'h00000000000000000000;
mem[5101] = 80'h00000000000000000000;
mem[5102] = 80'h10100000010000010010;
mem[5103] = 80'h00109400000208004500;
mem[5104] = 80'h0010002e2ac70000fffd;
mem[5105] = 80'h00100eb3c0550102c000;
mem[5106] = 80'h00100001ffabffabffab;
mem[5107] = 80'h00103857f87a50389aa0;
mem[5108] = 80'h0010d780f280cf482db2;
mem[5109] = 80'h0110dcc140960673862c;
mem[5110] = 80'h00000000000000000000;
mem[5111] = 80'h00000000000000000000;
mem[5112] = 80'h00000000000000000000;
mem[5113] = 80'h10100000010000010010;
mem[5114] = 80'h00109400000208004500;
mem[5115] = 80'h0010002e2ac80000fffd;
mem[5116] = 80'h00100eb2c0550102c000;
mem[5117] = 80'h00100001ffabffabffab;
mem[5118] = 80'h0010376faf832a68471e;
mem[5119] = 80'h00106d8c57b5435a9228;
mem[5120] = 80'h01100a96022c61b604e2;
mem[5121] = 80'h00000000000000000000;
mem[5122] = 80'h10100000010000010010;
mem[5123] = 80'h00109400000208004500;
mem[5124] = 80'h0010002e2ac90000fffd;
mem[5125] = 80'h00100eb1c0550102c000;
mem[5126] = 80'h00100001ffabffabffab;
mem[5127] = 80'h0010361e71aff21185a1;
mem[5128] = 80'h0010a65ed058b68ac879;
mem[5129] = 80'h01109a28509a75a08232;
mem[5130] = 80'h00000000000000000000;
mem[5131] = 80'h00000000000000000000;
mem[5132] = 80'h00000000000000000000;
mem[5133] = 80'h10100000010000010010;
mem[5134] = 80'h00109400000208004500;
mem[5135] = 80'h0010002e2aca0000fffd;
mem[5136] = 80'h00100eb0c0550102c000;
mem[5137] = 80'h00100001ffabffabffab;
mem[5138] = 80'h0010358c13da9a9bc261;
mem[5139] = 80'h0010fa29586ea8fb8d8b;
mem[5140] = 80'h0110dd5ef31d4112c0cc;
mem[5141] = 80'h00000000000000000000;
mem[5142] = 80'h00000000000000000000;
mem[5143] = 80'h00000000000000000000;
mem[5144] = 80'h10100000010000010010;
mem[5145] = 80'h00109400000208004500;
mem[5146] = 80'h0010002e2acb0000fffd;
mem[5147] = 80'h00100eafc0550102c000;
mem[5148] = 80'h00100001ffabffabffab;
mem[5149] = 80'h001034fdcdf642e200de;
mem[5150] = 80'h001031fbdf835d2bcbda;
mem[5151] = 80'h01100bfe72c8fc5f1eb3;
mem[5152] = 80'h00000000000000000000;
mem[5153] = 80'h10100000010000010010;
mem[5154] = 80'h00109400000208004500;
mem[5155] = 80'h0010002e2acc0000fffd;
mem[5156] = 80'h00100eaec0550102c000;
mem[5157] = 80'h00100001ffabffabffab;
mem[5158] = 80'h001033d9091c93f68f5e;
mem[5159] = 80'h00108914ceef61ca8f3f;
mem[5160] = 80'h01108fa9c6fd1ce307a8;
mem[5161] = 80'h00000000000000000000;
mem[5162] = 80'h00000000000000000000;
mem[5163] = 80'h00000000000000000000;
mem[5164] = 80'h00000000000000000000;
mem[5165] = 80'h10100000010000010010;
mem[5166] = 80'h00109400000208004500;
mem[5167] = 80'h0010002e2acd0000fffd;
mem[5168] = 80'h00100eadc0550102c000;
mem[5169] = 80'h00100001ffabffabffab;
mem[5170] = 80'h001032a8d7304b8f4de1;
mem[5171] = 80'h001042c64902941a8c6e;
mem[5172] = 80'h0110ab30053469f2f254;
mem[5173] = 80'h00000000000000000000;
mem[5174] = 80'h10100000010000010010;
mem[5175] = 80'h00109400000208004500;
mem[5176] = 80'h0010002e2ace0000fffd;
mem[5177] = 80'h00100eacc0550102c000;
mem[5178] = 80'h00100001ffabffabffab;
mem[5179] = 80'h0010313ab54523050a21;
mem[5180] = 80'h00101eb1c1348a6a0f9c;
mem[5181] = 80'h011067840ae95b8e09ea;
mem[5182] = 80'h00000000000000000000;
mem[5183] = 80'h00000000000000000000;
mem[5184] = 80'h00000000000000000000;
mem[5185] = 80'h00000000000000000000;
mem[5186] = 80'h10100000010000010010;
mem[5187] = 80'h00109400000208004500;
mem[5188] = 80'h0010002e2acf0000fffd;
mem[5189] = 80'h00100eabc0550102c000;
mem[5190] = 80'h00100001ffabffabffab;
mem[5191] = 80'h0010304b6b69fb7cc89e;
mem[5192] = 80'h0010d56346d97fba90cd;
mem[5193] = 80'h01101e9b54cf47a147dc;
mem[5194] = 80'h00000000000000000000;
mem[5195] = 80'h00000000000000000000;
mem[5196] = 80'h00000000000000000000;
mem[5197] = 80'h10100000010000010010;
mem[5198] = 80'h00109400000208004500;
mem[5199] = 80'h0010002e2ad00000fffd;
mem[5200] = 80'h00100eaac0550102c000;
mem[5201] = 80'h00100001ffabffabffab;
mem[5202] = 80'h00102f4a1ab7d7a4b15c;
mem[5203] = 80'h00106aa88b5f924f64a8;
mem[5204] = 80'h011014bc2b41e20c35d6;
mem[5205] = 80'h00000000000000000000;
mem[5206] = 80'h10100000010000010010;
mem[5207] = 80'h00109400000208004500;
mem[5208] = 80'h0010002e2ad10000fffd;
mem[5209] = 80'h00100ea9c0550102c000;
mem[5210] = 80'h00100001ffabffabffab;
mem[5211] = 80'h00102e3bc49b0fdd73e3;
mem[5212] = 80'h0010a17a0cb2679f6ff9;
mem[5213] = 80'h0110b98c4a168c60ed0b;
mem[5214] = 80'h00000000000000000000;
mem[5215] = 80'h00000000000000000000;
mem[5216] = 80'h00000000000000000000;
mem[5217] = 80'h10100000010000010010;
mem[5218] = 80'h00109400000208004500;
mem[5219] = 80'h0010002e2ad20000fffd;
mem[5220] = 80'h00100ea8c0550102c000;
mem[5221] = 80'h00100001ffabffabffab;
mem[5222] = 80'h00102da9a6ee67573423;
mem[5223] = 80'h0010fd0d848479efe50b;
mem[5224] = 80'h0110cfa0dfbee3ed17b8;
mem[5225] = 80'h00000000000000000000;
mem[5226] = 80'h00000000000000000000;
mem[5227] = 80'h00000000000000000000;
mem[5228] = 80'h10100000010000010010;
mem[5229] = 80'h00109400000208004500;
mem[5230] = 80'h0010002e2ad30000fffd;
mem[5231] = 80'h00100ea7c0550102c000;
mem[5232] = 80'h00100001ffabffabffab;
mem[5233] = 80'h00102cd878c2bf2ef69c;
mem[5234] = 80'h001036df03698c3f9b5a;
mem[5235] = 80'h0110953cad7a2ee6c5bf;
mem[5236] = 80'h00000000000000000000;
mem[5237] = 80'h10100000010000010010;
mem[5238] = 80'h00109400000208004500;
mem[5239] = 80'h0010002e2ad40000fffd;
mem[5240] = 80'h00100ea6c0550102c000;
mem[5241] = 80'h00100001ffabffabffab;
mem[5242] = 80'h00102bfcbc286e3a791c;
mem[5243] = 80'h00108e301205b0d929bf;
mem[5244] = 80'h01102d9c881992f39442;
mem[5245] = 80'h00000000000000000000;
mem[5246] = 80'h00000000000000000000;
mem[5247] = 80'h00000000000000000000;
mem[5248] = 80'h00000000000000000000;
mem[5249] = 80'h10100000010000010010;
mem[5250] = 80'h00109400000208004500;
mem[5251] = 80'h0010002e2ad50000fffd;
mem[5252] = 80'h00100ea5c0550102c000;
mem[5253] = 80'h00100001ffabffabffab;
mem[5254] = 80'h00102a8d6204b643bba3;
mem[5255] = 80'h001045e295e845096aee;
mem[5256] = 80'h011004c970fb0a49e84b;
mem[5257] = 80'h00000000000000000000;
mem[5258] = 80'h00000000000000000000;
mem[5259] = 80'h00000000000000000000;
mem[5260] = 80'h10100000010000010010;
mem[5261] = 80'h00109400000208004500;
mem[5262] = 80'h0010002e2ad60000fffd;
mem[5263] = 80'h00100ea4c0550102c000;
mem[5264] = 80'h00100001ffabffabffab;
mem[5265] = 80'h0010291f0071dec9fc63;
mem[5266] = 80'h001019951dde5b79b91c;
mem[5267] = 80'h0110c6c2e87542ef221b;
mem[5268] = 80'h00000000000000000000;
mem[5269] = 80'h00000000000000000000;
mem[5270] = 80'h00000000000000000000;
mem[5271] = 80'h10100000010000010010;
mem[5272] = 80'h00109400000208004500;
mem[5273] = 80'h0010002e2ad70000fffd;
mem[5274] = 80'h00100ea3c0550102c000;
mem[5275] = 80'h00100001ffabffabffab;
mem[5276] = 80'h0010286ede5d06b03edc;
mem[5277] = 80'h0010d2479a33aea9f84d;
mem[5278] = 80'h011089f5163fbe9c450c;
mem[5279] = 80'h00000000000000000000;
mem[5280] = 80'h10100000010000010010;
mem[5281] = 80'h00109400000208004500;
mem[5282] = 80'h0010002e2ad80000fffd;
mem[5283] = 80'h00100ea2c0550102c000;
mem[5284] = 80'h00100001ffabffabffab;
mem[5285] = 80'h0010275689a47ce0e362;
mem[5286] = 80'h0010684b3f0622bbc8d7;
mem[5287] = 80'h0110540407d94f4a9ed4;
mem[5288] = 80'h00000000000000000000;
mem[5289] = 80'h00000000000000000000;
mem[5290] = 80'h00000000000000000000;
mem[5291] = 80'h00000000000000000000;
mem[5292] = 80'h10100000010000010010;
mem[5293] = 80'h00109400000208004500;
mem[5294] = 80'h0010002e2ad90000fffd;
mem[5295] = 80'h00100ea1c0550102c000;
mem[5296] = 80'h00100001ffabffabffab;
mem[5297] = 80'h001026275788a49921dd;
mem[5298] = 80'h0010a399b8ebd76bb186;
mem[5299] = 80'h0110970f3f5248787758;
mem[5300] = 80'h00000000000000000000;
mem[5301] = 80'h10100000010000010010;
mem[5302] = 80'h00109400000208004500;
mem[5303] = 80'h0010002e2ada0000fffd;
mem[5304] = 80'h00100ea0c0550102c000;
mem[5305] = 80'h00100001ffabffabffab;
mem[5306] = 80'h001025b535fdcc13661d;
mem[5307] = 80'h0010ffee30ddc91b3874;
mem[5308] = 80'h0110b4708b4f10baa4c8;
mem[5309] = 80'h00000000000000000000;
mem[5310] = 80'h00000000000000000000;
mem[5311] = 80'h00000000000000000000;
mem[5312] = 80'h10100000010000010010;
mem[5313] = 80'h00109400000208004500;
mem[5314] = 80'h0010002e2adb0000fffd;
mem[5315] = 80'h00100e9fc0550102c000;
mem[5316] = 80'h00100001ffabffabffab;
mem[5317] = 80'h001024c4ebd1146aa4a2;
mem[5318] = 80'h0010343cb7303ccb3125;
mem[5319] = 80'h01107f225ddddef0f1df;
mem[5320] = 80'h00000000000000000000;
mem[5321] = 80'h00000000000000000000;
mem[5322] = 80'h00000000000000000000;
mem[5323] = 80'h10100000010000010010;
mem[5324] = 80'h00109400000208004500;
mem[5325] = 80'h0010002e2adc0000fffd;
mem[5326] = 80'h00100e9ec0550102c000;
mem[5327] = 80'h00100001ffabffabffab;
mem[5328] = 80'h001023e02f3bc57e2b22;
mem[5329] = 80'h00108cd3a65c002a54c0;
mem[5330] = 80'h0110cea26586932a177a;
mem[5331] = 80'h00000000000000000000;
mem[5332] = 80'h00000000000000000000;
mem[5333] = 80'h00000000000000000000;
mem[5334] = 80'h10100000010000010010;
mem[5335] = 80'h00109400000208004500;
mem[5336] = 80'h0010002e2add0000fffd;
mem[5337] = 80'h00100e9dc0550102c000;
mem[5338] = 80'h00100001ffabffabffab;
mem[5339] = 80'h00102291f1171d07e99d;
mem[5340] = 80'h0010470121b1f5fbd691;
mem[5341] = 80'h0110f5a2bace72dd0973;
mem[5342] = 80'h00000000000000000000;
mem[5343] = 80'h00000000000000000000;
mem[5344] = 80'h00000000000000000000;
mem[5345] = 80'h10100000010000010010;
mem[5346] = 80'h00109400000208004500;
mem[5347] = 80'h0010002e2ade0000fffd;
mem[5348] = 80'h00100e9cc0550102c000;
mem[5349] = 80'h00100001ffabffabffab;
mem[5350] = 80'h001021039362758dae5d;
mem[5351] = 80'h00101b76a987eb8b5463;
mem[5352] = 80'h01100a27189bbb635339;
mem[5353] = 80'h00000000000000000000;
mem[5354] = 80'h10100000010000010010;
mem[5355] = 80'h00109400000208004500;
mem[5356] = 80'h0010002e2adf0000fffd;
mem[5357] = 80'h00100e9bc0550102c000;
mem[5358] = 80'h00100001ffabffabffab;
mem[5359] = 80'h001020724d4eadf46ce2;
mem[5360] = 80'h0010d0a42e6a1e5b2a32;
mem[5361] = 80'h011050bbdf108fcf158b;
mem[5362] = 80'h00000000000000000000;
mem[5363] = 80'h00000000000000000000;
mem[5364] = 80'h00000000000000000000;
mem[5365] = 80'h10100000010000010010;
mem[5366] = 80'h00109400000208004500;
mem[5367] = 80'h0010002e2ae00000fffd;
mem[5368] = 80'h00100e9ac0550102c000;
mem[5369] = 80'h00100001ffabffabffab;
mem[5370] = 80'h00101f0170de2c3d5dd8;
mem[5371] = 80'h001064e1328a306089a9;
mem[5372] = 80'h0110e409b08b27e33871;
mem[5373] = 80'h00000000000000000000;
mem[5374] = 80'h00000000000000000000;
mem[5375] = 80'h00000000000000000000;
mem[5376] = 80'h10100000010000010010;
mem[5377] = 80'h00109400000208004500;
mem[5378] = 80'h0010002e2ae10000fffd;
mem[5379] = 80'h00100e99c0550102c000;
mem[5380] = 80'h00100001ffabffabffab;
mem[5381] = 80'h00101e70aef2f4449f67;
mem[5382] = 80'h0010af33b567c5b0c0f8;
mem[5383] = 80'h011022979114c12177b4;
mem[5384] = 80'h00000000000000000000;
mem[5385] = 80'h10100000010000010010;
mem[5386] = 80'h00109400000208004500;
mem[5387] = 80'h0010002e2ae20000fffd;
mem[5388] = 80'h00100e98c0550102c000;
mem[5389] = 80'h00100001ffabffabffab;
mem[5390] = 80'h00101de2cc879cced8a7;
mem[5391] = 80'h0010f3443d51dbc0950a;
mem[5392] = 80'h011051a2ad1b725bbbf7;
mem[5393] = 80'h00000000000000000000;
mem[5394] = 80'h00000000000000000000;
mem[5395] = 80'h00000000000000000000;
mem[5396] = 80'h00000000000000000000;
mem[5397] = 80'h00000000000000000000;
mem[5398] = 80'h10100000010000010010;
mem[5399] = 80'h00109400000208004500;
mem[5400] = 80'h0010002e2ae30000fffd;
mem[5401] = 80'h00100e97c0550102c000;
mem[5402] = 80'h00100001ffabffabffab;
mem[5403] = 80'h00101c9312ab44b71a18;
mem[5404] = 80'h00103896babc2e10d45b;
mem[5405] = 80'h01101e955d9e247bc1bf;
mem[5406] = 80'h00000000000000000000;
mem[5407] = 80'h10100000010000010010;
mem[5408] = 80'h00109400000208004500;
mem[5409] = 80'h0010002e2ae40000fffd;
mem[5410] = 80'h00100e96c0550102c000;
mem[5411] = 80'h00100001ffabffabffab;
mem[5412] = 80'h00101bb7d64195a39598;
mem[5413] = 80'h00108079abd012f1e7be;
mem[5414] = 80'h01100b0cb0c4e25d469a;
mem[5415] = 80'h00000000000000000000;
mem[5416] = 80'h00000000000000000000;
mem[5417] = 80'h00000000000000000000;
mem[5418] = 80'h10100000010000010010;
mem[5419] = 80'h00109400000208004500;
mem[5420] = 80'h0010002e2ae50000fffd;
mem[5421] = 80'h00100e95c0550102c000;
mem[5422] = 80'h00100001ffabffabffab;
mem[5423] = 80'h00101ac6086d4dda5727;
mem[5424] = 80'h00104bab2c3de721a4ef;
mem[5425] = 80'h011022591178947d9074;
mem[5426] = 80'h00000000000000000000;
mem[5427] = 80'h00000000000000000000;
mem[5428] = 80'h00000000000000000000;
mem[5429] = 80'h10100000010000010010;
mem[5430] = 80'h00109400000208004500;
mem[5431] = 80'h0010002e2ae60000fffd;
mem[5432] = 80'h00100e94c0550102c000;
mem[5433] = 80'h00100001ffabffabffab;
mem[5434] = 80'h001019546a18255010e7;
mem[5435] = 80'h001017dca40bf951161d;
mem[5436] = 80'h0110d849a2bbb85b03bc;
mem[5437] = 80'h00000000000000000000;
mem[5438] = 80'h00000000000000000000;
mem[5439] = 80'h00000000000000000000;
mem[5440] = 80'h10100000010000010010;
mem[5441] = 80'h00109400000208004500;
mem[5442] = 80'h0010002e2ae70000fffd;
mem[5443] = 80'h00100e93c0550102c000;
mem[5444] = 80'h00100001ffabffabffab;
mem[5445] = 80'h00101825b434fd29d258;
mem[5446] = 80'h0010dc0e23e60c82984c;
mem[5447] = 80'h0110c844f71ad8bf8bba;
mem[5448] = 80'h00000000000000000000;
mem[5449] = 80'h10100000010000010010;
mem[5450] = 80'h00109400000208004500;
mem[5451] = 80'h0010002e2ae80000fffd;
mem[5452] = 80'h00100e92c0550102c000;
mem[5453] = 80'h00100001ffabffabffab;
mem[5454] = 80'h0010171de3cd87790fe6;
mem[5455] = 80'h0010660286d3809067d6;
mem[5456] = 80'h011013df84999048d688;
mem[5457] = 80'h00000000000000000000;
mem[5458] = 80'h00000000000000000000;
mem[5459] = 80'h00000000000000000000;
mem[5460] = 80'h10100000010000010010;
mem[5461] = 80'h00109400000208004500;
mem[5462] = 80'h0010002e2ae90000fffd;
mem[5463] = 80'h00100e91c0550102c000;
mem[5464] = 80'h00100001ffabffabffab;
mem[5465] = 80'h0010166c3de15f00cd59;
mem[5466] = 80'h0010add0013e75407c87;
mem[5467] = 80'h0110bd9c20e5c985eb08;
mem[5468] = 80'h00000000000000000000;
mem[5469] = 80'h00000000000000000000;
mem[5470] = 80'h00000000000000000000;
mem[5471] = 80'h10100000010000010010;
mem[5472] = 80'h00109400000208004500;
mem[5473] = 80'h0010002e2aea0000fffd;
mem[5474] = 80'h00100e90c0550102c000;
mem[5475] = 80'h00100001ffabffabffab;
mem[5476] = 80'h001015fe5f94378a8a99;
mem[5477] = 80'h0010f1a789086b30f775;
mem[5478] = 80'h0110f881f27038962a50;
mem[5479] = 80'h00000000000000000000;
mem[5480] = 80'h00000000000000000000;
mem[5481] = 80'h00000000000000000000;
mem[5482] = 80'h10100000010000010010;
mem[5483] = 80'h00109400000208004500;
mem[5484] = 80'h0010002e2aeb0000fffd;
mem[5485] = 80'h00100e8fc0550102c000;
mem[5486] = 80'h00100001ffabffabffab;
mem[5487] = 80'h0010148f81b8eff34826;
mem[5488] = 80'h00103a750ee59ee07824;
mem[5489] = 80'h011082ed4e51db232356;
mem[5490] = 80'h00000000000000000000;
mem[5491] = 80'h10100000010000010010;
mem[5492] = 80'h00109400000208004500;
mem[5493] = 80'h0010002e2aec0000fffd;
mem[5494] = 80'h00100e8ec0550102c000;
mem[5495] = 80'h00100001ffabffabffab;
mem[5496] = 80'h001013ab45523ee7c7a6;
mem[5497] = 80'h0010829a1f89a2013bc1;
mem[5498] = 80'h01109f2d8160fccb8da3;
mem[5499] = 80'h00000000000000000000;
mem[5500] = 80'h00000000000000000000;
mem[5501] = 80'h00000000000000000000;
mem[5502] = 80'h10100000010000010010;
mem[5503] = 80'h00109400000208004500;
mem[5504] = 80'h0010002e2aed0000fffd;
mem[5505] = 80'h00100e8dc0550102c000;
mem[5506] = 80'h00100001ffabffabffab;
mem[5507] = 80'h001012da9b7ee69e0519;
mem[5508] = 80'h00104948986457d17890;
mem[5509] = 80'h0110b678fd67dc3a7e25;
mem[5510] = 80'h00000000000000000000;
mem[5511] = 80'h00000000000000000000;
mem[5512] = 80'h00000000000000000000;
mem[5513] = 80'h10100000010000010010;
mem[5514] = 80'h00109400000208004500;
mem[5515] = 80'h0010002e2aee0000fffd;
mem[5516] = 80'h00100e8cc0550102c000;
mem[5517] = 80'h00100001ffabffabffab;
mem[5518] = 80'h00101148f90b8e1442d9;
mem[5519] = 80'h0010153f105249a1bb62;
mem[5520] = 80'h011077008328a44127d6;
mem[5521] = 80'h00000000000000000000;
mem[5522] = 80'h00000000000000000000;
mem[5523] = 80'h00000000000000000000;
mem[5524] = 80'h10100000010000010010;
mem[5525] = 80'h00109400000208004500;
mem[5526] = 80'h0010002e2aef0000fffd;
mem[5527] = 80'h00100e8bc0550102c000;
mem[5528] = 80'h00100001ffabffabffab;
mem[5529] = 80'h001010392727566d8066;
mem[5530] = 80'h0010deed97bfbc71fa33;
mem[5531] = 80'h011038378c41d693806e;
mem[5532] = 80'h00000000000000000000;
mem[5533] = 80'h10100000010000010010;
mem[5534] = 80'h00109400000208004500;
mem[5535] = 80'h0010002e2af00000fffd;
mem[5536] = 80'h00100e8ac0550102c000;
mem[5537] = 80'h00100001ffabffabffab;
mem[5538] = 80'h00100f3856f97ab5f9a4;
mem[5539] = 80'h001061265a395185d056;
mem[5540] = 80'h011033081530d2661e65;
mem[5541] = 80'h00000000000000000000;
mem[5542] = 80'h00000000000000000000;
mem[5543] = 80'h00000000000000000000;
mem[5544] = 80'h00000000000000000000;
mem[5545] = 80'h10100000010000010010;
mem[5546] = 80'h00109400000208004500;
mem[5547] = 80'h0010002e2af10000fffd;
mem[5548] = 80'h00100e89c0550102c000;
mem[5549] = 80'h00100001ffabffabffab;
mem[5550] = 80'h00100e4988d5a2cc3b1b;
mem[5551] = 80'h0010aaf4ddd4a4559a07;
mem[5552] = 80'h0110a0c5230db1ffb789;
mem[5553] = 80'h00000000000000000000;
mem[5554] = 80'h00000000000000000000;
mem[5555] = 80'h00000000000000000000;
mem[5556] = 80'h10100000010000010010;
mem[5557] = 80'h00109400000208004500;
mem[5558] = 80'h0010002e2af20000fffd;
mem[5559] = 80'h00100e88c0550102c000;
mem[5560] = 80'h00100001ffabffabffab;
mem[5561] = 80'h00100ddbeaa0ca467cdb;
mem[5562] = 80'h0010f68355e2ba2550f5;
mem[5563] = 80'h0110db258dba862d70ee;
mem[5564] = 80'h00000000000000000000;
mem[5565] = 80'h10100000010000010010;
mem[5566] = 80'h00109400000208004500;
mem[5567] = 80'h0010002e2af30000fffd;
mem[5568] = 80'h00100e87c0550102c000;
mem[5569] = 80'h00100001ffabffabffab;
mem[5570] = 80'h00100caa348c123fbe64;
mem[5571] = 80'h00103d51d20f4ff52ea4;
mem[5572] = 80'h011081b9de71392e82f5;
mem[5573] = 80'h00000000000000000000;
mem[5574] = 80'h00000000000000000000;
mem[5575] = 80'h00000000000000000000;
mem[5576] = 80'h10100000010000010010;
mem[5577] = 80'h00109400000208004500;
mem[5578] = 80'h0010002e2af40000fffd;
mem[5579] = 80'h00100e86c0550102c000;
mem[5580] = 80'h00100001ffabffabffab;
mem[5581] = 80'h00100b8ef066c32b31e4;
mem[5582] = 80'h001085bec36373145f41;
mem[5583] = 80'h0110ff8ef3f3582ea6ee;
mem[5584] = 80'h00000000000000000000;
mem[5585] = 80'h00000000000000000000;
mem[5586] = 80'h00000000000000000000;
mem[5587] = 80'h10100000010000010010;
mem[5588] = 80'h00109400000208004500;
mem[5589] = 80'h0010002e2af50000fffd;
mem[5590] = 80'h00100e85c0550102c000;
mem[5591] = 80'h00100001ffabffabffab;
mem[5592] = 80'h00100aff2e4a1b52f35b;
mem[5593] = 80'h00104e6c448e86c4de10;
mem[5594] = 80'h0110a6ed194bf8da6903;
mem[5595] = 80'h00000000000000000000;
mem[5596] = 80'h00000000000000000000;
mem[5597] = 80'h00000000000000000000;
mem[5598] = 80'h10100000010000010010;
mem[5599] = 80'h00109400000208004500;
mem[5600] = 80'h0010002e2af60000fffd;
mem[5601] = 80'h00100e84c0550102c000;
mem[5602] = 80'h00100001ffabffabffab;
mem[5603] = 80'h0010096d4c3f73d8b49b;
mem[5604] = 80'h0010121bccb898b44be2;
mem[5605] = 80'h0110c38cfae7521bf506;
mem[5606] = 80'h00000000000000000000;
mem[5607] = 80'h10100000010000010010;
mem[5608] = 80'h00109400000208004500;
mem[5609] = 80'h0010002e2af70000fffd;
mem[5610] = 80'h00100e83c0550102c000;
mem[5611] = 80'h00100001ffabffabffab;
mem[5612] = 80'h0010081c9213aba17624;
mem[5613] = 80'h0010d9c94b556d6442b3;
mem[5614] = 80'h011008de65f5284be8c7;
mem[5615] = 80'h00000000000000000000;
mem[5616] = 80'h00000000000000000000;
mem[5617] = 80'h00000000000000000000;
mem[5618] = 80'h10100000010000010010;
mem[5619] = 80'h00109400000208004500;
mem[5620] = 80'h0010002e2af80000fffd;
mem[5621] = 80'h00100e82c0550102c000;
mem[5622] = 80'h00100001ffabffabffab;
mem[5623] = 80'h00100724c5ead1f1ab9a;
mem[5624] = 80'h001063c5ee60e176be29;
mem[5625] = 80'h011086163d87549ec25d;
mem[5626] = 80'h00000000000000000000;
mem[5627] = 80'h00000000000000000000;
mem[5628] = 80'h00000000000000000000;
mem[5629] = 80'h10100000010000010010;
mem[5630] = 80'h00109400000208004500;
mem[5631] = 80'h0010002e2af90000fffd;
mem[5632] = 80'h00100e81c0550102c000;
mem[5633] = 80'h00100001ffabffabffab;
mem[5634] = 80'h001006551bc609886925;
mem[5635] = 80'h0010a817698d14a6c678;
mem[5636] = 80'h0110762c08474b41e089;
mem[5637] = 80'h00000000000000000000;
mem[5638] = 80'h00000000000000000000;
mem[5639] = 80'h00000000000000000000;
mem[5640] = 80'h10100000010000010010;
mem[5641] = 80'h00109400000208004500;
mem[5642] = 80'h0010002e2afa0000fffd;
mem[5643] = 80'h00100e80c0550102c000;
mem[5644] = 80'h00100001ffabffabffab;
mem[5645] = 80'h001005c779b361022ee5;
mem[5646] = 80'h0010f460e1bb0ad9828a;
mem[5647] = 80'h0110196a73b35756c12d;
mem[5648] = 80'h00000000000000000000;
mem[5649] = 80'h10100000010000010010;
mem[5650] = 80'h00109400000208004500;
mem[5651] = 80'h0010002e2afb0000fffd;
mem[5652] = 80'h00100e7fc0550102c000;
mem[5653] = 80'h00100001ffabffabffab;
mem[5654] = 80'h001004b6a79fb97bec5a;
mem[5655] = 80'h00103fb26656ff09c3db;
mem[5656] = 80'h0110565dee87da13592f;
mem[5657] = 80'h00000000000000000000;
mem[5658] = 80'h00000000000000000000;
mem[5659] = 80'h00000000000000000000;
mem[5660] = 80'h00000000000000000000;
mem[5661] = 80'h10100000010000010010;
mem[5662] = 80'h00109400000208004500;
mem[5663] = 80'h0010002e2afc0000fffd;
mem[5664] = 80'h00100e7ec0550102c000;
mem[5665] = 80'h00100001ffabffabffab;
mem[5666] = 80'h001003926375686f63da;
mem[5667] = 80'h0010875d773ac3e8e13e;
mem[5668] = 80'h01107386b568100bf548;
mem[5669] = 80'h00000000000000000000;
mem[5670] = 80'h00000000000000000000;
mem[5671] = 80'h00000000000000000000;
mem[5672] = 80'h10100000010000010010;
mem[5673] = 80'h00109400000208004500;
mem[5674] = 80'h0010002e2afd0000fffd;
mem[5675] = 80'h00100e7dc0550102c000;
mem[5676] = 80'h00100001ffabffabffab;
mem[5677] = 80'h001002e3bd59b016a165;
mem[5678] = 80'h00104c8ff0d73638a36f;
mem[5679] = 80'h011069e26d5522510ace;
mem[5680] = 80'h00000000000000000000;
mem[5681] = 80'h10100000010000010010;
mem[5682] = 80'h00109400000208004500;
mem[5683] = 80'h0010002e2afe0000fffd;
mem[5684] = 80'h00100e7cc0550102c000;
mem[5685] = 80'h00100001ffabffabffab;
mem[5686] = 80'h00100171df2cd89ce6a5;
mem[5687] = 80'h001010f878e12848e19d;
mem[5688] = 80'h011080334c2c1bd809a9;
mem[5689] = 80'h00000000000000000000;
mem[5690] = 80'h00000000000000000000;
mem[5691] = 80'h00000000000000000000;
mem[5692] = 80'h10100000010000010010;
mem[5693] = 80'h00109400000208004500;
mem[5694] = 80'h0010002e2aff0000fffd;
mem[5695] = 80'h00100e7bc0550102c000;
mem[5696] = 80'h00100001ffabffabffab;
mem[5697] = 80'h00100000010000e5241a;
mem[5698] = 80'h0010db2aff0cdd989ecc;
mem[5699] = 80'h0110e99e99c4533f6bbb;
mem[5700] = 80'h00000000000000000000;
mem[5701] = 80'h00000000000000000000;
mem[5702] = 80'h00000000000000000000;
mem[5703] = 80'h10100000010000010010;
mem[5704] = 80'h00109400000208004500;
mem[5705] = 80'h0010002e2b000000fffd;
mem[5706] = 80'h00100e7ac0550102c000;
mem[5707] = 80'h00100001ffabffabffab;
mem[5708] = 80'h0010ff2f4b1bb732658f;
mem[5709] = 80'h00109d9a82578ed76603;
mem[5710] = 80'h011080af0376dd5c23c4;
mem[5711] = 80'h00000000000000000000;
mem[5712] = 80'h00000000000000000000;
mem[5713] = 80'h00000000000000000000;
mem[5714] = 80'h10100000010000010010;
mem[5715] = 80'h00109400000208004500;
mem[5716] = 80'h0010002e2b010000fffd;
mem[5717] = 80'h00100e79c0550102c000;
mem[5718] = 80'h00100001ffabffabffab;
mem[5719] = 80'h0010fe5e95376f4ba730;
mem[5720] = 80'h0010564805ba7b076d52;
mem[5721] = 80'h01102d9fe3f16d4bb0bd;
mem[5722] = 80'h00000000000000000000;
mem[5723] = 80'h10100000010000010010;
mem[5724] = 80'h00109400000208004500;
mem[5725] = 80'h0010002e2b020000fffd;
mem[5726] = 80'h00100e78c0550102c000;
mem[5727] = 80'h00100001ffabffabffab;
mem[5728] = 80'h0010fdccf74207c1e0f0;
mem[5729] = 80'h00100a3f8d8c6577e6a0;
mem[5730] = 80'h01106882d5d7428c0b8d;
mem[5731] = 80'h00000000000000000000;
mem[5732] = 80'h00000000000000000000;
mem[5733] = 80'h00000000000000000000;
mem[5734] = 80'h10100000010000010010;
mem[5735] = 80'h00109400000208004500;
mem[5736] = 80'h0010002e2b030000fffd;
mem[5737] = 80'h00100e77c0550102c000;
mem[5738] = 80'h00100001ffabffabffab;
mem[5739] = 80'h0010fcbd296edfb8224f;
mem[5740] = 80'h0010c1ed0a6190a679f1;
mem[5741] = 80'h011026adda37f727474f;
mem[5742] = 80'h00000000000000000000;
mem[5743] = 80'h00000000000000000000;
mem[5744] = 80'h00000000000000000000;
mem[5745] = 80'h10100000010000010010;
mem[5746] = 80'h00109400000208004500;
mem[5747] = 80'h0010002e2b040000fffd;
mem[5748] = 80'h00100e76c0550102c000;
mem[5749] = 80'h00100001ffabffabffab;
mem[5750] = 80'h0010fb99ed840eacadcf;
mem[5751] = 80'h001079021b0dac470914;
mem[5752] = 80'h01106baba54e9938eafa;
mem[5753] = 80'h00000000000000000000;
mem[5754] = 80'h00000000000000000000;
mem[5755] = 80'h00000000000000000000;
mem[5756] = 80'h10100000010000010010;
mem[5757] = 80'h00109400000208004500;
mem[5758] = 80'h0010002e2b050000fffd;
mem[5759] = 80'h00100e75c0550102c000;
mem[5760] = 80'h00100001ffabffabffab;
mem[5761] = 80'h0010fae833a8d6d56f70;
mem[5762] = 80'h0010b2d09ce059970945;
mem[5763] = 80'h01101a61be39a7e59a77;
mem[5764] = 80'h00000000000000000000;
mem[5765] = 80'h10100000010000010010;
mem[5766] = 80'h00109400000208004500;
mem[5767] = 80'h0010002e2b060000fffd;
mem[5768] = 80'h00100e74c0550102c000;
mem[5769] = 80'h00100001ffabffabffab;
mem[5770] = 80'h0010f97a51ddbe5f28b0;
mem[5771] = 80'h0010eea714d647e7bdb7;
mem[5772] = 80'h01104ad779a387ad97cf;
mem[5773] = 80'h00000000000000000000;
mem[5774] = 80'h00000000000000000000;
mem[5775] = 80'h00000000000000000000;
mem[5776] = 80'h00000000000000000000;
mem[5777] = 80'h10100000010000010010;
mem[5778] = 80'h00109400000208004500;
mem[5779] = 80'h0010002e2b070000fffd;
mem[5780] = 80'h00100e73c0550102c000;
mem[5781] = 80'h00100001ffabffabffab;
mem[5782] = 80'h0010f80b8ff16626ea0f;
mem[5783] = 80'h00102575933bb237f4e6;
mem[5784] = 80'h01108c493bb3169a95b1;
mem[5785] = 80'h00000000000000000000;
mem[5786] = 80'h00000000000000000000;
mem[5787] = 80'h00000000000000000000;
mem[5788] = 80'h10100000010000010010;
mem[5789] = 80'h00109400000208004500;
mem[5790] = 80'h0010002e2b080000fffd;
mem[5791] = 80'h00100e72c0550102c000;
mem[5792] = 80'h00100001ffabffabffab;
mem[5793] = 80'h0010f733d8081c7637b1;
mem[5794] = 80'h00109f79360e3e25cb7c;
mem[5795] = 80'h01104186bbebe74477a2;
mem[5796] = 80'h00000000000000000000;
mem[5797] = 80'h10100000010000010010;
mem[5798] = 80'h00109400000208004500;
mem[5799] = 80'h0010002e2b090000fffd;
mem[5800] = 80'h00100e71c0550102c000;
mem[5801] = 80'h00100001ffabffabffab;
mem[5802] = 80'h0010f6420624c40ff50e;
mem[5803] = 80'h001054abb1e3cbf5912d;
mem[5804] = 80'h0110d138158fba4f25a2;
mem[5805] = 80'h00000000000000000000;
mem[5806] = 80'h00000000000000000000;
mem[5807] = 80'h00000000000000000000;
mem[5808] = 80'h10100000010000010010;
mem[5809] = 80'h00109400000208004500;
mem[5810] = 80'h0010002e2b0a0000fffd;
mem[5811] = 80'h00100e70c0550102c000;
mem[5812] = 80'h00100001ffabffabffab;
mem[5813] = 80'h0010f5d06451ac85b2ce;
mem[5814] = 80'h001008dc39d5d58554df;
mem[5815] = 80'h0110bae61e8c648f2455;
mem[5816] = 80'h00000000000000000000;
mem[5817] = 80'h10100000010000010010;
mem[5818] = 80'h00109400000208004500;
mem[5819] = 80'h0010002e2b0b0000fffd;
mem[5820] = 80'h00100e6fc0550102c000;
mem[5821] = 80'h00100001ffabffabffab;
mem[5822] = 80'h0010f4a1ba7d74fc7071;
mem[5823] = 80'h0010c30ebe382055158e;
mem[5824] = 80'h0110f5d1be753a8bacb1;
mem[5825] = 80'h00000000000000000000;
mem[5826] = 80'h00000000000000000000;
mem[5827] = 80'h00000000000000000000;
mem[5828] = 80'h00000000000000000000;
mem[5829] = 80'h10100000010000010010;
mem[5830] = 80'h00109400000208004500;
mem[5831] = 80'h0010002e2b0c0000fffd;
mem[5832] = 80'h00100e6ec0550102c000;
mem[5833] = 80'h00100001ffabffabffab;
mem[5834] = 80'h0010f3857e97a5e8fff1;
mem[5835] = 80'h00107be1af541cb4546b;
mem[5836] = 80'h01108e73bd3ee7754b8b;
mem[5837] = 80'h00000000000000000000;
mem[5838] = 80'h00000000000000000000;
mem[5839] = 80'h00000000000000000000;
mem[5840] = 80'h10100000010000010010;
mem[5841] = 80'h00109400000208004500;
mem[5842] = 80'h0010002e2b0d0000fffd;
mem[5843] = 80'h00100e6dc0550102c000;
mem[5844] = 80'h00100001ffabffabffab;
mem[5845] = 80'h0010f2f4a0bb7d913d4e;
mem[5846] = 80'h0010b03328b9e967d53a;
mem[5847] = 80'h01108e408b9f91d733c4;
mem[5848] = 80'h00000000000000000000;
mem[5849] = 80'h00000000000000000000;
mem[5850] = 80'h00000000000000000000;
mem[5851] = 80'h10100000010000010010;
mem[5852] = 80'h00109400000208004500;
mem[5853] = 80'h0010002e2b0e0000fffd;
mem[5854] = 80'h00100e6cc0550102c000;
mem[5855] = 80'h00100001ffabffabffab;
mem[5856] = 80'h0010f166c2ce151b7a8e;
mem[5857] = 80'h0010ec44a08ff71750c8;
mem[5858] = 80'h0110e852ff18da88c714;
mem[5859] = 80'h00000000000000000000;
mem[5860] = 80'h10100000010000010010;
mem[5861] = 80'h00109400000208004500;
mem[5862] = 80'h0010002e2b0f0000fffd;
mem[5863] = 80'h00100e6bc0550102c000;
mem[5864] = 80'h00100001ffabffabffab;
mem[5865] = 80'h0010f0171ce2cd62b831;
mem[5866] = 80'h00102796276202c74899;
mem[5867] = 80'h01101342bfd6beefa017;
mem[5868] = 80'h00000000000000000000;
mem[5869] = 80'h00000000000000000000;
mem[5870] = 80'h00000000000000000000;
mem[5871] = 80'h10100000010000010010;
mem[5872] = 80'h00109400000208004500;
mem[5873] = 80'h0010002e2b100000fffd;
mem[5874] = 80'h00100e6ac0550102c000;
mem[5875] = 80'h00100001ffabffabffab;
mem[5876] = 80'h0010ef166d3ce1bac1f3;
mem[5877] = 80'h0010985deae4ef32bffc;
mem[5878] = 80'h01104c368155355dbc9e;
mem[5879] = 80'h00000000000000000000;
mem[5880] = 80'h10100000010000010010;
mem[5881] = 80'h00109400000208004500;
mem[5882] = 80'h0010002e2b110000fffd;
mem[5883] = 80'h00100e69c0550102c000;
mem[5884] = 80'h00100001ffabffabffab;
mem[5885] = 80'h0010ee67b31039c3034c;
mem[5886] = 80'h0010538f6d091ae237ad;
mem[5887] = 80'h0110afcd5e8294018faa;
mem[5888] = 80'h00000000000000000000;
mem[5889] = 80'h00000000000000000000;
mem[5890] = 80'h00000000000000000000;
mem[5891] = 80'h00000000000000000000;
mem[5892] = 80'h10100000010000010010;
mem[5893] = 80'h00109400000208004500;
mem[5894] = 80'h0010002e2b120000fffd;
mem[5895] = 80'h00100e68c0550102c000;
mem[5896] = 80'h00100001ffabffabffab;
mem[5897] = 80'h0010edf5d1655149448c;
mem[5898] = 80'h00100ff8e53f0492bc5f;
mem[5899] = 80'h0110ead009d461edd7b6;
mem[5900] = 80'h00000000000000000000;
mem[5901] = 80'h00000000000000000000;
mem[5902] = 80'h00000000000000000000;
mem[5903] = 80'h10100000010000010010;
mem[5904] = 80'h00109400000208004500;
mem[5905] = 80'h0010002e2b130000fffd;
mem[5906] = 80'h00100e67c0550102c000;
mem[5907] = 80'h00100001ffabffabffab;
mem[5908] = 80'h0010ec840f4989308633;
mem[5909] = 80'h0010c42a62d2f142c20e;
mem[5910] = 80'h0110b04c6a325884bc37;
mem[5911] = 80'h00000000000000000000;
mem[5912] = 80'h00000000000000000000;
mem[5913] = 80'h00000000000000000000;
mem[5914] = 80'h10100000010000010010;
mem[5915] = 80'h00109400000208004500;
mem[5916] = 80'h0010002e2b140000fffd;
mem[5917] = 80'h00100e66c0550102c000;
mem[5918] = 80'h00100001ffabffabffab;
mem[5919] = 80'h0010eba0cba3582409b3;
mem[5920] = 80'h00107cc573becda3f0eb;
mem[5921] = 80'h011096e4a0eb2cc924b0;
mem[5922] = 80'h00000000000000000000;
mem[5923] = 80'h10100000010000010010;
mem[5924] = 80'h00109400000208004500;
mem[5925] = 80'h0010002e2b150000fffd;
mem[5926] = 80'h00100e65c0550102c000;
mem[5927] = 80'h00100001ffabffabffab;
mem[5928] = 80'h0010ead1158f805dcb0c;
mem[5929] = 80'h0010b717f4533873b3ba;
mem[5930] = 80'h0110bfb15ce9c8543e7d;
mem[5931] = 80'h00000000000000000000;
mem[5932] = 80'h00000000000000000000;
mem[5933] = 80'h00000000000000000000;
mem[5934] = 80'h10100000010000010010;
mem[5935] = 80'h00109400000208004500;
mem[5936] = 80'h0010002e2b160000fffd;
mem[5937] = 80'h00100e64c0550102c000;
mem[5938] = 80'h00100001ffabffabffab;
mem[5939] = 80'h0010e94377fae8d78ccc;
mem[5940] = 80'h0010eb607c652602e048;
mem[5941] = 80'h0110511269f9558da2a4;
mem[5942] = 80'h00000000000000000000;
mem[5943] = 80'h00000000000000000000;
mem[5944] = 80'h00000000000000000000;
mem[5945] = 80'h10100000010000010010;
mem[5946] = 80'h00109400000208004500;
mem[5947] = 80'h0010002e2b170000fffd;
mem[5948] = 80'h00100e63c0550102c000;
mem[5949] = 80'h00100001ffabffabffab;
mem[5950] = 80'h0010e832a9d630ae4e73;
mem[5951] = 80'h001020b2fb88d3d2af19;
mem[5952] = 80'h01103d2a128396843950;
mem[5953] = 80'h00000000000000000000;
mem[5954] = 80'h00000000000000000000;
mem[5955] = 80'h00000000000000000000;
mem[5956] = 80'h10100000010000010010;
mem[5957] = 80'h00109400000208004500;
mem[5958] = 80'h0010002e2b180000fffd;
mem[5959] = 80'h00100e62c0550102c000;
mem[5960] = 80'h00100001ffabffabffab;
mem[5961] = 80'h0010e70afe2f4afe93cd;
mem[5962] = 80'h00109abe5ebd5fc01183;
mem[5963] = 80'h0110d84cf8ec065ab702;
mem[5964] = 80'h00000000000000000000;
mem[5965] = 80'h00000000000000000000;
mem[5966] = 80'h00000000000000000000;
mem[5967] = 80'h10100000010000010010;
mem[5968] = 80'h00109400000208004500;
mem[5969] = 80'h0010002e2b190000fffd;
mem[5970] = 80'h00100e61c0550102c000;
mem[5971] = 80'h00100001ffabffabffab;
mem[5972] = 80'h0010e67b200392875172;
mem[5973] = 80'h0010516cd950aa106ad2;
mem[5974] = 80'h01107d2558c15478a510;
mem[5975] = 80'h00000000000000000000;
mem[5976] = 80'h10100000010000010010;
mem[5977] = 80'h00109400000208004500;
mem[5978] = 80'h0010002e2b1a0000fffd;
mem[5979] = 80'h00100e60c0550102c000;
mem[5980] = 80'h00100001ffabffabffab;
mem[5981] = 80'h0010e5e94276fa0d16b2;
mem[5982] = 80'h00100d1b5166b460ee20;
mem[5983] = 80'h011028069dd6ef20ebc1;
mem[5984] = 80'h00000000000000000000;
mem[5985] = 80'h00000000000000000000;
mem[5986] = 80'h00000000000000000000;
mem[5987] = 80'h10100000010000010010;
mem[5988] = 80'h00109400000208004500;
mem[5989] = 80'h0010002e2b1b0000fffd;
mem[5990] = 80'h00100e5fc0550102c000;
mem[5991] = 80'h00100001ffabffabffab;
mem[5992] = 80'h0010e4989c5a2274d40d;
mem[5993] = 80'h0010c6c9d68b41b06e71;
mem[5994] = 80'h01104254f8be28b75688;
mem[5995] = 80'h00000000000000000000;
mem[5996] = 80'h10100000010000010010;
mem[5997] = 80'h00109400000208004500;
mem[5998] = 80'h0010002e2b1c0000fffd;
mem[5999] = 80'h00100e5ec0550102c000;
mem[6000] = 80'h00100001ffabffabffab;
mem[6001] = 80'h0010e3bc58b0f3605b8d;
mem[6002] = 80'h00107e26c7e77d510e94;
mem[6003] = 80'h01100c21968f8839f151;
mem[6004] = 80'h00000000000000000000;
mem[6005] = 80'h00000000000000000000;
mem[6006] = 80'h00000000000000000000;
mem[6007] = 80'h10100000010000010010;
mem[6008] = 80'h00109400000208004500;
mem[6009] = 80'h0010002e2b1d0000fffd;
mem[6010] = 80'h00100e5dc0550102c000;
mem[6011] = 80'h00100001ffabffabffab;
mem[6012] = 80'h0010e2cd869c2b199932;
mem[6013] = 80'h0010b5f4400a888101c5;
mem[6014] = 80'h01106dd5e42e696eb488;
mem[6015] = 80'h00000000000000000000;
mem[6016] = 80'h00000000000000000000;
mem[6017] = 80'h00000000000000000000;
mem[6018] = 80'h10100000010000010010;
mem[6019] = 80'h00109400000208004500;
mem[6020] = 80'h0010002e2b1e0000fffd;
mem[6021] = 80'h00100e5cc0550102c000;
mem[6022] = 80'h00100001ffabffabffab;
mem[6023] = 80'h0010e15fe4e94393def2;
mem[6024] = 80'h0010e983c83c96f18d37;
mem[6025] = 80'h0110b15f8fe6c375b9d5;
mem[6026] = 80'h00000000000000000000;
mem[6027] = 80'h00000000000000000000;
mem[6028] = 80'h00000000000000000000;
mem[6029] = 80'h10100000010000010010;
mem[6030] = 80'h00109400000208004500;
mem[6031] = 80'h0010002e2b1f0000fffd;
mem[6032] = 80'h00100e5bc0550102c000;
mem[6033] = 80'h00100001ffabffabffab;
mem[6034] = 80'h0010e02e3ac59bea1c4d;
mem[6035] = 80'h001022514fd16321f366;
mem[6036] = 80'h0110ebc37865366762b6;
mem[6037] = 80'h00000000000000000000;
mem[6038] = 80'h00000000000000000000;
mem[6039] = 80'h00000000000000000000;
mem[6040] = 80'h10100000010000010010;
mem[6041] = 80'h00109400000208004500;
mem[6042] = 80'h0010002e2b200000fffd;
mem[6043] = 80'h00100e5ac0550102c000;
mem[6044] = 80'h00100001ffabffabffab;
mem[6045] = 80'h0010df5d07551a232d77;
mem[6046] = 80'h0010961453314d1dd0fd;
mem[6047] = 80'h0110c17908d8842d83db;
mem[6048] = 80'h00000000000000000000;
mem[6049] = 80'h10100000010000010010;
mem[6050] = 80'h00109400000208004500;
mem[6051] = 80'h0010002e2b210000fffd;
mem[6052] = 80'h00100e59c0550102c000;
mem[6053] = 80'h00100001ffabffabffab;
mem[6054] = 80'h0010de2cd979c25aefc8;
mem[6055] = 80'h00105dc6d4dcb8cd99ac;
mem[6056] = 80'h011007e70931c91f2e32;
mem[6057] = 80'h00000000000000000000;
mem[6058] = 80'h00000000000000000000;
mem[6059] = 80'h00000000000000000000;
mem[6060] = 80'h00000000000000000000;
mem[6061] = 80'h10100000010000010010;
mem[6062] = 80'h00109400000208004500;
mem[6063] = 80'h0010002e2b220000fffd;
mem[6064] = 80'h00100e58c0550102c000;
mem[6065] = 80'h00100001ffabffabffab;
mem[6066] = 80'h0010ddbebb0caad0a808;
mem[6067] = 80'h001001b15ceaa6bd4c5e;
mem[6068] = 80'h01106f4a5359ae703bfb;
mem[6069] = 80'h00000000000000000000;
mem[6070] = 80'h00000000000000000000;
mem[6071] = 80'h00000000000000000000;
mem[6072] = 80'h10100000010000010010;
mem[6073] = 80'h00109400000208004500;
mem[6074] = 80'h0010002e2b230000fffd;
mem[6075] = 80'h00100e57c0550102c000;
mem[6076] = 80'h00100001ffabffabffab;
mem[6077] = 80'h0010dccf652072a96ab7;
mem[6078] = 80'h0010ca63db07536d0d0f;
mem[6079] = 80'h0110207dba492b9e24a8;
mem[6080] = 80'h00000000000000000000;
mem[6081] = 80'h10100000010000010010;
mem[6082] = 80'h00109400000208004500;
mem[6083] = 80'h0010002e2b240000fffd;
mem[6084] = 80'h00100e56c0550102c000;
mem[6085] = 80'h00100001ffabffabffab;
mem[6086] = 80'h0010dbeba1caa3bde537;
mem[6087] = 80'h0010728cca6b6f8cbcea;
mem[6088] = 80'h0110481e47c673b7a643;
mem[6089] = 80'h00000000000000000000;
mem[6090] = 80'h00000000000000000000;
mem[6091] = 80'h00000000000000000000;
mem[6092] = 80'h10100000010000010010;
mem[6093] = 80'h00109400000208004500;
mem[6094] = 80'h0010002e2b250000fffd;
mem[6095] = 80'h00100e55c0550102c000;
mem[6096] = 80'h00100001ffabffabffab;
mem[6097] = 80'h0010da9a7fe67bc42788;
mem[6098] = 80'h0010b95e4d869a5cfcbb;
mem[6099] = 80'h01103418301c262c7eca;
mem[6100] = 80'h00000000000000000000;
mem[6101] = 80'h00000000000000000000;
mem[6102] = 80'h00000000000000000000;
mem[6103] = 80'h10100000010000010010;
mem[6104] = 80'h00109400000208004500;
mem[6105] = 80'h0010002e2b260000fffd;
mem[6106] = 80'h00100e54c0550102c000;
mem[6107] = 80'h00100001ffabffabffab;
mem[6108] = 80'h0010d9081d93134e6048;
mem[6109] = 80'h0010e529c5b0842c4849;
mem[6110] = 80'h011064aeb9ce2fcf8e64;
mem[6111] = 80'h00000000000000000000;
mem[6112] = 80'h10100000010000010010;
mem[6113] = 80'h00109400000208004500;
mem[6114] = 80'h0010002e2b270000fffd;
mem[6115] = 80'h00100e53c0550102c000;
mem[6116] = 80'h00100001ffabffabffab;
mem[6117] = 80'h0010d879c3bfcb37a2f7;
mem[6118] = 80'h00102efb425d71fc4018;
mem[6119] = 80'h01109ccd355caa56af25;
mem[6120] = 80'h00000000000000000000;
mem[6121] = 80'h00000000000000000000;
mem[6122] = 80'h00000000000000000000;
mem[6123] = 80'h00000000000000000000;
mem[6124] = 80'h10100000010000010010;
mem[6125] = 80'h00109400000208004500;
mem[6126] = 80'h0010002e2b280000fffd;
mem[6127] = 80'h00100e52c0550102c000;
mem[6128] = 80'h00100001ffabffabffab;
mem[6129] = 80'h0010d7419446b1677f49;
mem[6130] = 80'h001094f7e768fdeebc82;
mem[6131] = 80'h011012051aefc19e9833;
mem[6132] = 80'h00000000000000000000;
mem[6133] = 80'h10100000010000010010;
mem[6134] = 80'h00109400000208004500;
mem[6135] = 80'h0010002e2b290000fffd;
mem[6136] = 80'h00100e51c0550102c000;
mem[6137] = 80'h00100001ffabffabffab;
mem[6138] = 80'h0010d6304a6a691ebdf6;
mem[6139] = 80'h00105f256085083f25d3;
mem[6140] = 80'h0110f68cd4056cf345a8;
mem[6141] = 80'h00000000000000000000;
mem[6142] = 80'h00000000000000000000;
mem[6143] = 80'h00000000000000000000;
mem[6144] = 80'h00000000000000000000;
mem[6145] = 80'h10100000010000010010;
mem[6146] = 80'h00109400000208004500;
mem[6147] = 80'h0010002e2b2a0000fffd;
mem[6148] = 80'h00100e50c0550102c000;
mem[6149] = 80'h00100001ffabffabffab;
mem[6150] = 80'h0010d5a2281f0194fa36;
mem[6151] = 80'h00100352e8b3164fae21;
mem[6152] = 80'h0110b391a26a72828767;
mem[6153] = 80'h00000000000000000000;
mem[6154] = 80'h00000000000000000000;
mem[6155] = 80'h00000000000000000000;
mem[6156] = 80'h10100000010000010010;
mem[6157] = 80'h00109400000208004500;
mem[6158] = 80'h0010002e2b2b0000fffd;
mem[6159] = 80'h00100e4fc0550102c000;
mem[6160] = 80'h00100001ffabffabffab;
mem[6161] = 80'h0010d4d3f633d9ed3889;
mem[6162] = 80'h0010c8806f5ee39fa170;
mem[6163] = 80'h0110d265932bc19db9c8;
mem[6164] = 80'h00000000000000000000;
mem[6165] = 80'h10100000010000010010;
mem[6166] = 80'h00109400000208004500;
mem[6167] = 80'h0010002e2b2c0000fffd;
mem[6168] = 80'h00100e4ec0550102c000;
mem[6169] = 80'h00100001ffabffabffab;
mem[6170] = 80'h0010d3f732d908f9b709;
mem[6171] = 80'h0010706f7e32df7ee295;
mem[6172] = 80'h0110cfa5b8cf5565bcf1;
mem[6173] = 80'h00000000000000000000;
mem[6174] = 80'h00000000000000000000;
mem[6175] = 80'h00000000000000000000;
mem[6176] = 80'h00000000000000000000;
mem[6177] = 80'h10100000010000010010;
mem[6178] = 80'h00109400000208004500;
mem[6179] = 80'h0010002e2b2d0000fffd;
mem[6180] = 80'h00100e4dc0550102c000;
mem[6181] = 80'h00100001ffabffabffab;
mem[6182] = 80'h0010d286ecf5d08075b6;
mem[6183] = 80'h0010bbbdf9df2aaea1c4;
mem[6184] = 80'h0110e6f0914a68df35b3;
mem[6185] = 80'h00000000000000000000;
mem[6186] = 80'h00000000000000000000;
mem[6187] = 80'h00000000000000000000;
mem[6188] = 80'h10100000010000010010;
mem[6189] = 80'h00109400000208004500;
mem[6190] = 80'h0010002e2b2e0000fffd;
mem[6191] = 80'h00100e4cc0550102c000;
mem[6192] = 80'h00100001ffabffabffab;
mem[6193] = 80'h0010d1148e80b80a3276;
mem[6194] = 80'h0010e7ca71e934dee236;
mem[6195] = 80'h01103c1009109f393d4f;
mem[6196] = 80'h00000000000000000000;
mem[6197] = 80'h10100000010000010010;
mem[6198] = 80'h00109400000208004500;
mem[6199] = 80'h0010002e2b2f0000fffd;
mem[6200] = 80'h00100e4bc0550102c000;
mem[6201] = 80'h00100001ffabffabffab;
mem[6202] = 80'h0010d06550ac6073f0c9;
mem[6203] = 80'h00102c18f604c10ebd67;
mem[6204] = 80'h0110535b99c1671bfc00;
mem[6205] = 80'h00000000000000000000;
mem[6206] = 80'h00000000000000000000;
mem[6207] = 80'h00000000000000000000;
mem[6208] = 80'h00000000000000000000;
mem[6209] = 80'h10100000010000010010;
mem[6210] = 80'h00109400000208004500;
mem[6211] = 80'h0010002e2b300000fffd;
mem[6212] = 80'h00100e4ac0550102c000;
mem[6213] = 80'h00100001ffabffabffab;
mem[6214] = 80'h0010cf6421724cab890b;
mem[6215] = 80'h001093d33b822cfb0a02;
mem[6216] = 80'h011001e3313cde65c17c;
mem[6217] = 80'h00000000000000000000;
mem[6218] = 80'h10100000010000010010;
mem[6219] = 80'h00109400000208004500;
mem[6220] = 80'h0010002e2b310000fffd;
mem[6221] = 80'h00100e49c0550102c000;
mem[6222] = 80'h00100001ffabffabffab;
mem[6223] = 80'h0010ce15ff5e94d24bb4;
mem[6224] = 80'h00105801bc6fd92b4253;
mem[6225] = 80'h0110f44c2dc78a41d295;
mem[6226] = 80'h00000000000000000000;
mem[6227] = 80'h00000000000000000000;
mem[6228] = 80'h00000000000000000000;
mem[6229] = 80'h00000000000000000000;
mem[6230] = 80'h10100000010000010010;
mem[6231] = 80'h00109400000208004500;
mem[6232] = 80'h0010002e2b320000fffd;
mem[6233] = 80'h00100e48c0550102c000;
mem[6234] = 80'h00100001ffabffabffab;
mem[6235] = 80'h0010cd879d2bfc580c74;
mem[6236] = 80'h001004763459c75bf6a1;
mem[6237] = 80'h0110a4faf0b717f82ddd;
mem[6238] = 80'h00000000000000000000;
mem[6239] = 80'h10100000010000010010;
mem[6240] = 80'h00109400000208004500;
mem[6241] = 80'h0010002e2b330000fffd;
mem[6242] = 80'h00100e47c0550102c000;
mem[6243] = 80'h00100001ffabffabffab;
mem[6244] = 80'h0010ccf643072421cecb;
mem[6245] = 80'h0010cfa4b3b4328875f0;
mem[6246] = 80'h0110c2ab0e97ac50c051;
mem[6247] = 80'h00000000000000000000;
mem[6248] = 80'h00000000000000000000;
mem[6249] = 80'h00000000000000000000;
mem[6250] = 80'h00000000000000000000;
mem[6251] = 80'h10100000010000010010;
mem[6252] = 80'h00109400000208004500;
mem[6253] = 80'h0010002e2b340000fffd;
mem[6254] = 80'h00100e46c0550102c000;
mem[6255] = 80'h00100001ffabffabffab;
mem[6256] = 80'h0010cbd287edf535414b;
mem[6257] = 80'h0010774ba2d80e690615;
mem[6258] = 80'h0110dafe6c1daf9d082b;
mem[6259] = 80'h00000000000000000000;
mem[6260] = 80'h00000000000000000000;
mem[6261] = 80'h00000000000000000000;
mem[6262] = 80'h10100000010000010010;
mem[6263] = 80'h00109400000208004500;
mem[6264] = 80'h0010002e2b350000fffd;
mem[6265] = 80'h00100e45c0550102c000;
mem[6266] = 80'h00100001ffabffabffab;
mem[6267] = 80'h0010caa359c12d4c83f4;
mem[6268] = 80'h0010bc992535fbb91944;
mem[6269] = 80'h0110b8797b13a9907aeb;
mem[6270] = 80'h00000000000000000000;
mem[6271] = 80'h10100000010000010010;
mem[6272] = 80'h00109400000208004500;
mem[6273] = 80'h0010002e2b360000fffd;
mem[6274] = 80'h00100e44c0550102c000;
mem[6275] = 80'h00100001ffabffabffab;
mem[6276] = 80'h0010c9313bb445c6c434;
mem[6277] = 80'h0010e0eead03e5c992b6;
mem[6278] = 80'h0110fd64ed46e9cbcabc;
mem[6279] = 80'h00000000000000000000;
mem[6280] = 80'h00000000000000000000;
mem[6281] = 80'h00000000000000000000;
mem[6282] = 80'h00000000000000000000;
mem[6283] = 80'h10100000010000010010;
mem[6284] = 80'h00109400000208004500;
mem[6285] = 80'h0010002e2b370000fffd;
mem[6286] = 80'h00100e43c0550102c000;
mem[6287] = 80'h00100001ffabffabffab;
mem[6288] = 80'h0010c840e5989dbf068b;
mem[6289] = 80'h00102b3c2aee10191be7;
mem[6290] = 80'h01102daefe021b954102;
mem[6291] = 80'h00000000000000000000;
mem[6292] = 80'h00000000000000000000;
mem[6293] = 80'h00000000000000000000;
mem[6294] = 80'h10100000010000010010;
mem[6295] = 80'h00109400000208004500;
mem[6296] = 80'h0010002e2b380000fffd;
mem[6297] = 80'h00100e42c0550102c000;
mem[6298] = 80'h00100001ffabffabffab;
mem[6299] = 80'h0010c778b261e7efdb35;
mem[6300] = 80'h001091308fdb9c0be77d;
mem[6301] = 80'h0110a3667b03b3dbf165;
mem[6302] = 80'h00000000000000000000;
mem[6303] = 80'h10100000010000010010;
mem[6304] = 80'h00109400000208004500;
mem[6305] = 80'h0010002e2b390000fffd;
mem[6306] = 80'h00100e41c0550102c000;
mem[6307] = 80'h00100001ffabffabffab;
mem[6308] = 80'h0010c6096c4d3f96198a;
mem[6309] = 80'h00105ae2083669db9f2c;
mem[6310] = 80'h0110535cb50b587624d3;
mem[6311] = 80'h00000000000000000000;
mem[6312] = 80'h00000000000000000000;
mem[6313] = 80'h00000000000000000000;
mem[6314] = 80'h10100000010000010010;
mem[6315] = 80'h00109400000208004500;
mem[6316] = 80'h0010002e2b3a0000fffd;
mem[6317] = 80'h00100e40c0550102c000;
mem[6318] = 80'h00100001ffabffabffab;
mem[6319] = 80'h0010c59b0e38571c5e4a;
mem[6320] = 80'h00100695800077ab5bde;
mem[6321] = 80'h01100bb310f33807a532;
mem[6322] = 80'h00000000000000000000;
mem[6323] = 80'h00000000000000000000;
mem[6324] = 80'h00000000000000000000;
mem[6325] = 80'h10100000010000010010;
mem[6326] = 80'h00109400000208004500;
mem[6327] = 80'h0010002e2b3b0000fffd;
mem[6328] = 80'h00100e3fc0550102c000;
mem[6329] = 80'h00100001ffabffabffab;
mem[6330] = 80'h0010c4ead0148f659cf5;
mem[6331] = 80'h0010cd4707ed827b1b8f;
mem[6332] = 80'h011077b553b06d6dcdff;
mem[6333] = 80'h00000000000000000000;
mem[6334] = 80'h00000000000000000000;
mem[6335] = 80'h00000000000000000000;
mem[6336] = 80'h10100000010000010010;
mem[6337] = 80'h00109400000208004500;
mem[6338] = 80'h0010002e2b3c0000fffd;
mem[6339] = 80'h00100e3ec0550102c000;
mem[6340] = 80'h00100001ffabffabffab;
mem[6341] = 80'h0010c3ce14fe5e711375;
mem[6342] = 80'h001075a81681be9bba6a;
mem[6343] = 80'h01102b958487e3e6aa16;
mem[6344] = 80'h00000000000000000000;
mem[6345] = 80'h10100000010000010010;
mem[6346] = 80'h00109400000208004500;
mem[6347] = 80'h0010002e2b3d0000fffd;
mem[6348] = 80'h00100e3dc0550102c000;
mem[6349] = 80'h00100001ffabffabffab;
mem[6350] = 80'h0010c2bfcad28608d1ca;
mem[6351] = 80'h0010be7a916c4b4bfb3b;
mem[6352] = 80'h011064a21f89d6dc6ce0;
mem[6353] = 80'h00000000000000000000;
mem[6354] = 80'h00000000000000000000;
mem[6355] = 80'h00000000000000000000;
mem[6356] = 80'h10100000010000010010;
mem[6357] = 80'h00109400000208004500;
mem[6358] = 80'h0010002e2b3e0000fffd;
mem[6359] = 80'h00100e3cc0550102c000;
mem[6360] = 80'h00100001ffabffabffab;
mem[6361] = 80'h0010c12da8a7ee82960a;
mem[6362] = 80'h0010e20d195a553b3ec9;
mem[6363] = 80'h01100f7c72b482cdabe5;
mem[6364] = 80'h00000000000000000000;
mem[6365] = 80'h00000000000000000000;
mem[6366] = 80'h00000000000000000000;
mem[6367] = 80'h10100000010000010010;
mem[6368] = 80'h00109400000208004500;
mem[6369] = 80'h0010002e2b3f0000fffd;
mem[6370] = 80'h00100e3bc0550102c000;
mem[6371] = 80'h00100001ffabffabffab;
mem[6372] = 80'h0010c05c768b36fb54b5;
mem[6373] = 80'h001029df9eb7a0eb4798;
mem[6374] = 80'h0110cc77bfd42f82cbbf;
mem[6375] = 80'h00000000000000000000;
mem[6376] = 80'h00000000000000000000;
mem[6377] = 80'h00000000000000000000;
mem[6378] = 80'h10100000010000010010;
mem[6379] = 80'h00109400000208004500;
mem[6380] = 80'h0010002e2b400000fffd;
mem[6381] = 80'h00100e3ac0550102c000;
mem[6382] = 80'h00100001ffabffabffab;
mem[6383] = 80'h0010bfcbd386ed10f47f;
mem[6384] = 80'h00108a87209a094c8fff;
mem[6385] = 80'h0110cf5e7750ebb356f4;
mem[6386] = 80'h00000000000000000000;
mem[6387] = 80'h10100000010000010010;
mem[6388] = 80'h00109400000208004500;
mem[6389] = 80'h0010002e2b410000fffd;
mem[6390] = 80'h00100e39c0550102c000;
mem[6391] = 80'h00100001ffabffabffab;
mem[6392] = 80'h0010beba0daa356936c0;
mem[6393] = 80'h00104155a777fc9c06ae;
mem[6394] = 80'h01101f94bbc529853335;
mem[6395] = 80'h00000000000000000000;
mem[6396] = 80'h00000000000000000000;
mem[6397] = 80'h00000000000000000000;
mem[6398] = 80'h00000000000000000000;
mem[6399] = 80'h10100000010000010010;
mem[6400] = 80'h00109400000208004500;
mem[6401] = 80'h0010002e2b420000fffd;
mem[6402] = 80'h00100e38c0550102c000;
mem[6403] = 80'h00100001ffabffabffab;
mem[6404] = 80'h0010bd286fdf5de37100;
mem[6405] = 80'h00101d222f41e2ec8d5c;
mem[6406] = 80'h01105a89ecdd4b050fb8;
mem[6407] = 80'h00000000000000000000;
mem[6408] = 80'h00000000000000000000;
mem[6409] = 80'h00000000000000000000;
mem[6410] = 80'h10100000010000010010;
mem[6411] = 80'h00109400000208004500;
mem[6412] = 80'h0010002e2b430000fffd;
mem[6413] = 80'h00100e37c0550102c000;
mem[6414] = 80'h00100001ffabffabffab;
mem[6415] = 80'h0010bc59b1f3859ab3bf;
mem[6416] = 80'h0010d6f0a8ac173c920d;
mem[6417] = 80'h0110380ef762fc36712a;
mem[6418] = 80'h00000000000000000000;
mem[6419] = 80'h10100000010000010010;
mem[6420] = 80'h00109400000208004500;
mem[6421] = 80'h0010002e2b440000fffd;
mem[6422] = 80'h00100e36c0550102c000;
mem[6423] = 80'h00100001ffabffabffab;
mem[6424] = 80'h0010bb7d7519548e3c3f;
mem[6425] = 80'h00106e1fb9c02bdde2e8;
mem[6426] = 80'h0110750892ecf6b4280c;
mem[6427] = 80'h00000000000000000000;
mem[6428] = 80'h00000000000000000000;
mem[6429] = 80'h00000000000000000000;
mem[6430] = 80'h10100000010000010010;
mem[6431] = 80'h00109400000208004500;
mem[6432] = 80'h0010002e2b450000fffd;
mem[6433] = 80'h00100e35c0550102c000;
mem[6434] = 80'h00100001ffabffabffab;
mem[6435] = 80'h0010ba0cab358cf7fe80;
mem[6436] = 80'h0010a5cd3e2dde3262b9;
mem[6437] = 80'h0110f6cef38e74fabb5c;
mem[6438] = 80'h00000000000000000000;
mem[6439] = 80'h10100000010000010010;
mem[6440] = 80'h00109400000208004500;
mem[6441] = 80'h0010002e2b460000fffd;
mem[6442] = 80'h00100e34c0550102c000;
mem[6443] = 80'h00100001ffabffabffab;
mem[6444] = 80'h0010b99ec940e47db940;
mem[6445] = 80'h0010f9bab61bc042d64b;
mem[6446] = 80'h0110a678f2837bc47d17;
mem[6447] = 80'h00000000000000000000;
mem[6448] = 80'h00000000000000000000;
mem[6449] = 80'h00000000000000000000;
mem[6450] = 80'h00000000000000000000;
mem[6451] = 80'h10100000010000010010;
mem[6452] = 80'h00109400000208004500;
mem[6453] = 80'h0010002e2b470000fffd;
mem[6454] = 80'h00100e33c0550102c000;
mem[6455] = 80'h00100001ffabffabffab;
mem[6456] = 80'h0010b8ef176c3c047bff;
mem[6457] = 80'h0010326831f635929d1a;
mem[6458] = 80'h011006843a11bd7773b3;
mem[6459] = 80'h00000000000000000000;
mem[6460] = 80'h00000000000000000000;
mem[6461] = 80'h00000000000000000000;
mem[6462] = 80'h10100000010000010010;
mem[6463] = 80'h00109400000208004500;
mem[6464] = 80'h0010002e2b480000fffd;
mem[6465] = 80'h00100e32c0550102c000;
mem[6466] = 80'h00100001ffabffabffab;
mem[6467] = 80'h0010b7d740954654a641;
mem[6468] = 80'h0010886494c3b9802380;
mem[6469] = 80'h0110e3e23cf17c8b316e;
mem[6470] = 80'h00000000000000000000;
mem[6471] = 80'h00000000000000000000;
mem[6472] = 80'h00000000000000000000;
mem[6473] = 80'h10100000010000010010;
mem[6474] = 80'h00109400000208004500;
mem[6475] = 80'h0010002e2b490000fffd;
mem[6476] = 80'h00100e31c0550102c000;
mem[6477] = 80'h00100001ffabffabffab;
mem[6478] = 80'h0010b6a69eb99e2d64fe;
mem[6479] = 80'h001043b6132e4c507cd1;
mem[6480] = 80'h01108ca9fac336b3887c;
mem[6481] = 80'h00000000000000000000;
mem[6482] = 80'h10100000010000010010;
mem[6483] = 80'h00109400000208004500;
mem[6484] = 80'h0010002e2b4a0000fffd;
mem[6485] = 80'h00100e30c0550102c000;
mem[6486] = 80'h00100001ffabffabffab;
mem[6487] = 80'h0010b534fcccf6a7233e;
mem[6488] = 80'h00101fc19b1852203f23;
mem[6489] = 80'h0110564991b1454fa48a;
mem[6490] = 80'h00000000000000000000;
mem[6491] = 80'h00000000000000000000;
mem[6492] = 80'h00000000000000000000;
mem[6493] = 80'h10100000010000010010;
mem[6494] = 80'h00109400000208004500;
mem[6495] = 80'h0010002e2b4b0000fffd;
mem[6496] = 80'h00100e2fc0550102c000;
mem[6497] = 80'h00100001ffabffabffab;
mem[6498] = 80'h0010b44522e02edee181;
mem[6499] = 80'h0010d4131cf5a7f07c72;
mem[6500] = 80'h01107f1c83f1939ab412;
mem[6501] = 80'h00000000000000000000;
mem[6502] = 80'h10100000010000010010;
mem[6503] = 80'h00109400000208004500;
mem[6504] = 80'h0010002e2b4c0000fffd;
mem[6505] = 80'h00100e2ec0550102c000;
mem[6506] = 80'h00100001ffabffabffab;
mem[6507] = 80'h0010b361e60affca6e01;
mem[6508] = 80'h00106cfc0d999b113e97;
mem[6509] = 80'h011051ed529b5ace89c3;
mem[6510] = 80'h00000000000000000000;
mem[6511] = 80'h00000000000000000000;
mem[6512] = 80'h00000000000000000000;
mem[6513] = 80'h00000000000000000000;
mem[6514] = 80'h10100000010000010010;
mem[6515] = 80'h00109400000208004500;
mem[6516] = 80'h0010002e2b4d0000fffd;
mem[6517] = 80'h00100e2dc0550102c000;
mem[6518] = 80'h00100001ffabffabffab;
mem[6519] = 80'h0010b210382627b3acbe;
mem[6520] = 80'h0010a72e8a746ec130c6;
mem[6521] = 80'h011003286d0415be1192;
mem[6522] = 80'h00000000000000000000;
mem[6523] = 80'h00000000000000000000;
mem[6524] = 80'h00000000000000000000;
mem[6525] = 80'h00000000000000000000;
mem[6526] = 80'h10100000010000010010;
mem[6527] = 80'h00109400000208004500;
mem[6528] = 80'h0010002e2b4e0000fffd;
mem[6529] = 80'h00100e2cc0550102c000;
mem[6530] = 80'h00100001ffabffabffab;
mem[6531] = 80'h0010b1825a534f39eb7e;
mem[6532] = 80'h0010fb59024270b1bb34;
mem[6533] = 80'h0110463549ba9f128a24;
mem[6534] = 80'h00000000000000000000;
mem[6535] = 80'h00000000000000000000;
mem[6536] = 80'h00000000000000000000;
mem[6537] = 80'h10100000010000010010;
mem[6538] = 80'h00109400000208004500;
mem[6539] = 80'h0010002e2b4f0000fffd;
mem[6540] = 80'h00100e2bc0550102c000;
mem[6541] = 80'h00100001ffabffabffab;
mem[6542] = 80'h0010b0f3847f974029c1;
mem[6543] = 80'h0010308b85af85602365;
mem[6544] = 80'h0110918d18fd5d6e1865;
mem[6545] = 80'h00000000000000000000;
mem[6546] = 80'h10100000010000010010;
mem[6547] = 80'h00109400000208004500;
mem[6548] = 80'h0010002e2b500000fffd;
mem[6549] = 80'h00100e2ac0550102c000;
mem[6550] = 80'h00100001ffabffabffab;
mem[6551] = 80'h0010aff2f5a1bb985003;
mem[6552] = 80'h00108f4048296895d400;
mem[6553] = 80'h0110cef96bd5fe97d7e8;
mem[6554] = 80'h00000000000000000000;
mem[6555] = 80'h00000000000000000000;
mem[6556] = 80'h00000000000000000000;
mem[6557] = 80'h10100000010000010010;
mem[6558] = 80'h00109400000208004500;
mem[6559] = 80'h0010002e2b510000fffd;
mem[6560] = 80'h00100e29c0550102c000;
mem[6561] = 80'h00100001ffabffabffab;
mem[6562] = 80'h0010ae832b8d63e192bc;
mem[6563] = 80'h00104492cfc49d45dc51;
mem[6564] = 80'h0110369a6ac86e2546d2;
mem[6565] = 80'h00000000000000000000;
mem[6566] = 80'h10100000010000010010;
mem[6567] = 80'h00109400000208004500;
mem[6568] = 80'h0010002e2b520000fffd;
mem[6569] = 80'h00100e28c0550102c000;
mem[6570] = 80'h00100001ffabffabffab;
mem[6571] = 80'h0010ad1149f80b6bd57c;
mem[6572] = 80'h001018e547f2833569a3;
mem[6573] = 80'h0110551d8540e1b9c4c8;
mem[6574] = 80'h00000000000000000000;
mem[6575] = 80'h00000000000000000000;
mem[6576] = 80'h00000000000000000000;
mem[6577] = 80'h10100000010000010010;
mem[6578] = 80'h00109400000208004500;
mem[6579] = 80'h0010002e2b530000fffd;
mem[6580] = 80'h00100e27c0550102c000;
mem[6581] = 80'h00100001ffabffabffab;
mem[6582] = 80'h0010ac6097d4d31217c3;
mem[6583] = 80'h0010d337c01f76e528f2;
mem[6584] = 80'h01101a2a839b7fa38b4e;
mem[6585] = 80'h00000000000000000000;
mem[6586] = 80'h00000000000000000000;
mem[6587] = 80'h00000000000000000000;
mem[6588] = 80'h10100000010000010010;
mem[6589] = 80'h00109400000208004500;
mem[6590] = 80'h0010002e2b540000fffd;
mem[6591] = 80'h00100e26c0550102c000;
mem[6592] = 80'h00100001ffabffabffab;
mem[6593] = 80'h0010ab44533e02069843;
mem[6594] = 80'h00106bd8d1734a049917;
mem[6595] = 80'h01107249d4818fb98471;
mem[6596] = 80'h00000000000000000000;
mem[6597] = 80'h00000000000000000000;
mem[6598] = 80'h00000000000000000000;
mem[6599] = 80'h10100000010000010010;
mem[6600] = 80'h00109400000208004500;
mem[6601] = 80'h0010002e2b550000fffd;
mem[6602] = 80'h00100e25c0550102c000;
mem[6603] = 80'h00100001ffabffabffab;
mem[6604] = 80'h0010aa358d12da7f5afc;
mem[6605] = 80'h0010a00a569ebfd4d846;
mem[6606] = 80'h01103d7ec6f8274462a3;
mem[6607] = 80'h00000000000000000000;
mem[6608] = 80'h10100000010000010010;
mem[6609] = 80'h00109400000208004500;
mem[6610] = 80'h0010002e2b560000fffd;
mem[6611] = 80'h00100e24c0550102c000;
mem[6612] = 80'h00100001ffabffabffab;
mem[6613] = 80'h0010a9a7ef67b2f51d3c;
mem[6614] = 80'h0010fc7ddea8a1a40db4;
mem[6615] = 80'h011055d3b66bfccc732f;
mem[6616] = 80'h00000000000000000000;
mem[6617] = 80'h00000000000000000000;
mem[6618] = 80'h00000000000000000000;
mem[6619] = 80'h00000000000000000000;
mem[6620] = 80'h10100000010000010010;
mem[6621] = 80'h00109400000208004500;
mem[6622] = 80'h0010002e2b570000fffd;
mem[6623] = 80'h00100e23c0550102c000;
mem[6624] = 80'h00100001ffabffabffab;
mem[6625] = 80'h0010a8d6314b6a8cdf83;
mem[6626] = 80'h001037af5945547447e5;
mem[6627] = 80'h0110c61ee8600b72de29;
mem[6628] = 80'h00000000000000000000;
mem[6629] = 80'h00000000000000000000;
mem[6630] = 80'h00000000000000000000;
mem[6631] = 80'h10100000010000010010;
mem[6632] = 80'h00109400000208004500;
mem[6633] = 80'h0010002e2b580000fffd;
mem[6634] = 80'h00100e22c0550102c000;
mem[6635] = 80'h00100001ffabffabffab;
mem[6636] = 80'h0010a7ee66b210dc023d;
mem[6637] = 80'h00108da3fc70d865787f;
mem[6638] = 80'h01105281b0cad8043fcb;
mem[6639] = 80'h00000000000000000000;
mem[6640] = 80'h10100000010000010010;
mem[6641] = 80'h00109400000208004500;
mem[6642] = 80'h0010002e2b590000fffd;
mem[6643] = 80'h00100e21c0550102c000;
mem[6644] = 80'h00100001ffabffabffab;
mem[6645] = 80'h0010a69fb89ec8a5c082;
mem[6646] = 80'h001046717b9d2db5062e;
mem[6647] = 80'h0110081d198a5fa62b06;
mem[6648] = 80'h00000000000000000000;
mem[6649] = 80'h00000000000000000000;
mem[6650] = 80'h00000000000000000000;
mem[6651] = 80'h00000000000000000000;
mem[6652] = 80'h10100000010000010010;
mem[6653] = 80'h00109400000208004500;
mem[6654] = 80'h0010002e2b5a0000fffd;
mem[6655] = 80'h00100e20c0550102c000;
mem[6656] = 80'h00100001ffabffabffab;
mem[6657] = 80'h0010a50ddaeba02f8742;
mem[6658] = 80'h00101a06f3ab33c585dc;
mem[6659] = 80'h0110c4a9cc96de05642f;
mem[6660] = 80'h00000000000000000000;
mem[6661] = 80'h00000000000000000000;
mem[6662] = 80'h00000000000000000000;
mem[6663] = 80'h10100000010000010010;
mem[6664] = 80'h00109400000208004500;
mem[6665] = 80'h0010002e2b5b0000fffd;
mem[6666] = 80'h00100e1fc0550102c000;
mem[6667] = 80'h00100001ffabffabffab;
mem[6668] = 80'h0010a47c04c7785645fd;
mem[6669] = 80'h0010d1d47446c615858d;
mem[6670] = 80'h0110b56351461cefae15;
mem[6671] = 80'h00000000000000000000;
mem[6672] = 80'h10100000010000010010;
mem[6673] = 80'h00109400000208004500;
mem[6674] = 80'h0010002e2b5c0000fffd;
mem[6675] = 80'h00100e1ec0550102c000;
mem[6676] = 80'h00100001ffabffabffab;
mem[6677] = 80'h0010a358c02da942ca7d;
mem[6678] = 80'h0010693b652afaf4e568;
mem[6679] = 80'h0110fb167edeb404618a;
mem[6680] = 80'h00000000000000000000;
mem[6681] = 80'h00000000000000000000;
mem[6682] = 80'h00000000000000000000;
mem[6683] = 80'h10100000010000010010;
mem[6684] = 80'h00109400000208004500;
mem[6685] = 80'h0010002e2b5d0000fffd;
mem[6686] = 80'h00100e1dc0550102c000;
mem[6687] = 80'h00100001ffabffabffab;
mem[6688] = 80'h0010a2291e01713b08c2;
mem[6689] = 80'h0010a2e9e2c70f246a39;
mem[6690] = 80'h0110817a454e2d8ae949;
mem[6691] = 80'h00000000000000000000;
mem[6692] = 80'h10100000010000010010;
mem[6693] = 80'h00109400000208004500;
mem[6694] = 80'h0010002e2b5e0000fffd;
mem[6695] = 80'h00100e1cc0550102c000;
mem[6696] = 80'h00100001ffabffabffab;
mem[6697] = 80'h0010a1bb7c7419b14f02;
mem[6698] = 80'h0010fe9e6af11154e1cb;
mem[6699] = 80'h0110c4675804189d264b;
mem[6700] = 80'h00000000000000000000;
mem[6701] = 80'h00000000000000000000;
mem[6702] = 80'h00000000000000000000;
mem[6703] = 80'h00000000000000000000;
mem[6704] = 80'h10100000010000010010;
mem[6705] = 80'h00109400000208004500;
mem[6706] = 80'h0010002e2b5f0000fffd;
mem[6707] = 80'h00100e1bc0550102c000;
mem[6708] = 80'h00100001ffabffabffab;
mem[6709] = 80'h0010a0caa258c1c88dbd;
mem[6710] = 80'h0010354ced1ce4849a9a;
mem[6711] = 80'h0110610e6abf0132b58b;
mem[6712] = 80'h00000000000000000000;
mem[6713] = 80'h00000000000000000000;
mem[6714] = 80'h00000000000000000000;
mem[6715] = 80'h10100000010000010010;
mem[6716] = 80'h00109400000208004500;
mem[6717] = 80'h0010002e2b600000fffd;
mem[6718] = 80'h00100e1ac0550102c000;
mem[6719] = 80'h00100001ffabffabffab;
mem[6720] = 80'h00109fb99fc84001bc87;
mem[6721] = 80'h00108109f1fccabf3b01;
mem[6722] = 80'h0110b3de974eed685e87;
mem[6723] = 80'h00000000000000000000;
mem[6724] = 80'h00000000000000000000;
mem[6725] = 80'h00000000000000000000;
mem[6726] = 80'h10100000010000010010;
mem[6727] = 80'h00109400000208004500;
mem[6728] = 80'h0010002e2b610000fffd;
mem[6729] = 80'h00100e19c0550102c000;
mem[6730] = 80'h00100001ffabffabffab;
mem[6731] = 80'h00109ec841e498787e38;
mem[6732] = 80'h00104adb76113f6f7450;
mem[6733] = 80'h0110dfe6b40e623c314f;
mem[6734] = 80'h00000000000000000000;
mem[6735] = 80'h10100000010000010010;
mem[6736] = 80'h00109400000208004500;
mem[6737] = 80'h0010002e2b620000fffd;
mem[6738] = 80'h00100e18c0550102c000;
mem[6739] = 80'h00100001ffabffabffab;
mem[6740] = 80'h00109d5a2391f0f239f8;
mem[6741] = 80'h001016acfe27211e26a2;
mem[6742] = 80'h01100274b520ee008de0;
mem[6743] = 80'h00000000000000000000;
mem[6744] = 80'h00000000000000000000;
mem[6745] = 80'h00000000000000000000;
mem[6746] = 80'h10100000010000010010;
mem[6747] = 80'h00109400000208004500;
mem[6748] = 80'h0010002e2b630000fffd;
mem[6749] = 80'h00100e17c0550102c000;
mem[6750] = 80'h00100001ffabffabffab;
mem[6751] = 80'h00109c2bfdbd288bfb47;
mem[6752] = 80'h0010dd7e79cad4ce64f3;
mem[6753] = 80'h01101810992770557192;
mem[6754] = 80'h00000000000000000000;
mem[6755] = 80'h00000000000000000000;
mem[6756] = 80'h00000000000000000000;
mem[6757] = 80'h10100000010000010010;
mem[6758] = 80'h00109400000208004500;
mem[6759] = 80'h0010002e2b640000fffd;
mem[6760] = 80'h00100e16c0550102c000;
mem[6761] = 80'h00100001ffabffabffab;
mem[6762] = 80'h00109b0f3957f99f74c7;
mem[6763] = 80'h0010659168a6e82f5616;
mem[6764] = 80'h01103eb871fbabaa31c2;
mem[6765] = 80'h00000000000000000000;
mem[6766] = 80'h00000000000000000000;
mem[6767] = 80'h00000000000000000000;
mem[6768] = 80'h10100000010000010010;
mem[6769] = 80'h00109400000208004500;
mem[6770] = 80'h0010002e2b650000fffd;
mem[6771] = 80'h00100e15c0550102c000;
mem[6772] = 80'h00100001ffabffabffab;
mem[6773] = 80'h00109a7ee77b21e6b678;
mem[6774] = 80'h0010ae43ef4b1dff2947;
mem[6775] = 80'h0110571569bb989c90fe;
mem[6776] = 80'h00000000000000000000;
mem[6777] = 80'h00000000000000000000;
mem[6778] = 80'h00000000000000000000;
mem[6779] = 80'h10100000010000010010;
mem[6780] = 80'h00109400000208004500;
mem[6781] = 80'h0010002e2b660000fffd;
mem[6782] = 80'h00100e14c0550102c000;
mem[6783] = 80'h00100001ffabffabffab;
mem[6784] = 80'h001099ec850e496cf1b8;
mem[6785] = 80'h0010f234677d038fa3b5;
mem[6786] = 80'h0110213983af698b1a27;
mem[6787] = 80'h00000000000000000000;
mem[6788] = 80'h10100000010000010010;
mem[6789] = 80'h00109400000208004500;
mem[6790] = 80'h0010002e2b670000fffd;
mem[6791] = 80'h00100e13c0550102c000;
mem[6792] = 80'h00100001ffabffabffab;
mem[6793] = 80'h0010989d5b2291153307;
mem[6794] = 80'h001039e6e090f65f2be4;
mem[6795] = 80'h0110c2c248a556fd7f4d;
mem[6796] = 80'h00000000000000000000;
mem[6797] = 80'h00000000000000000000;
mem[6798] = 80'h00000000000000000000;
mem[6799] = 80'h10100000010000010010;
mem[6800] = 80'h00109400000208004500;
mem[6801] = 80'h0010002e2b680000fffd;
mem[6802] = 80'h00100e12c0550102c000;
mem[6803] = 80'h00100001ffabffabffab;
mem[6804] = 80'h001097a50cdbeb45eeb9;
mem[6805] = 80'h001083ea45a57a4dd77e;
mem[6806] = 80'h01104c0a1a19172f6651;
mem[6807] = 80'h00000000000000000000;
mem[6808] = 80'h00000000000000000000;
mem[6809] = 80'h00000000000000000000;
mem[6810] = 80'h10100000010000010010;
mem[6811] = 80'h00109400000208004500;
mem[6812] = 80'h0010002e2b690000fffd;
mem[6813] = 80'h00100e11c0550102c000;
mem[6814] = 80'h00100001ffabffabffab;
mem[6815] = 80'h001096d4d2f7333c2c06;
mem[6816] = 80'h00104838c2488f9dce2f;
mem[6817] = 80'h0110842b4a7725a1e44a;
mem[6818] = 80'h00000000000000000000;
mem[6819] = 80'h00000000000000000000;
mem[6820] = 80'h00000000000000000000;
mem[6821] = 80'h10100000010000010010;
mem[6822] = 80'h00109400000208004500;
mem[6823] = 80'h0010002e2b6a0000fffd;
mem[6824] = 80'h00100e10c0550102c000;
mem[6825] = 80'h00100001ffabffabffab;
mem[6826] = 80'h00109546b0825bb66bc6;
mem[6827] = 80'h0010144f4a7e91ed4bdd;
mem[6828] = 80'h0110e239d3e708f613f2;
mem[6829] = 80'h00000000000000000000;
mem[6830] = 80'h10100000010000010010;
mem[6831] = 80'h00109400000208004500;
mem[6832] = 80'h0010002e2b6b0000fffd;
mem[6833] = 80'h00100e0fc0550102c000;
mem[6834] = 80'h00100001ffabffabffab;
mem[6835] = 80'h001094376eae83cfa979;
mem[6836] = 80'h0010df9dcd93643aca8c;
mem[6837] = 80'h01103ecab50dac9399e2;
mem[6838] = 80'h00000000000000000000;
mem[6839] = 80'h00000000000000000000;
mem[6840] = 80'h00000000000000000000;
mem[6841] = 80'h10100000010000010010;
mem[6842] = 80'h00109400000208004500;
mem[6843] = 80'h0010002e2b6c0000fffd;
mem[6844] = 80'h00100e0ec0550102c000;
mem[6845] = 80'h00100001ffabffabffab;
mem[6846] = 80'h00109313aa4452db26f9;
mem[6847] = 80'h00106772dcff58db8b69;
mem[6848] = 80'h01104568dab3494fe1dc;
mem[6849] = 80'h00000000000000000000;
mem[6850] = 80'h00000000000000000000;
mem[6851] = 80'h00000000000000000000;
mem[6852] = 80'h10100000010000010010;
mem[6853] = 80'h00109400000208004500;
mem[6854] = 80'h0010002e2b6d0000fffd;
mem[6855] = 80'h00100e0dc0550102c000;
mem[6856] = 80'h00100001ffabffabffab;
mem[6857] = 80'h0010926274688aa2e446;
mem[6858] = 80'h0010aca05b12ad0bc538;
mem[6859] = 80'h01101a61f5f2116f57c3;
mem[6860] = 80'h00000000000000000000;
mem[6861] = 80'h00000000000000000000;
mem[6862] = 80'h00000000000000000000;
mem[6863] = 80'h10100000010000010010;
mem[6864] = 80'h00109400000208004500;
mem[6865] = 80'h0010002e2b6e0000fffd;
mem[6866] = 80'h00100e0cc0550102c000;
mem[6867] = 80'h00100001ffabffabffab;
mem[6868] = 80'h001091f0161de228a386;
mem[6869] = 80'h0010f0d7d324b37b0fca;
mem[6870] = 80'h01106181e97e389868c3;
mem[6871] = 80'h00000000000000000000;
mem[6872] = 80'h10100000010000010010;
mem[6873] = 80'h00109400000208004500;
mem[6874] = 80'h0010002e2b6f0000fffd;
mem[6875] = 80'h00100e0bc0550102c000;
mem[6876] = 80'h00100001ffabffabffab;
mem[6877] = 80'h00109081c8313a516139;
mem[6878] = 80'h00103b0554c946ab559b;
mem[6879] = 80'h0110f13fee6c6e13038d;
mem[6880] = 80'h00000000000000000000;
mem[6881] = 80'h00000000000000000000;
mem[6882] = 80'h00000000000000000000;
mem[6883] = 80'h10100000010000010010;
mem[6884] = 80'h00109400000208004500;
mem[6885] = 80'h0010002e2b700000fffd;
mem[6886] = 80'h00100e0ac0550102c000;
mem[6887] = 80'h00100001ffabffabffab;
mem[6888] = 80'h00108f80b9ef168918fb;
mem[6889] = 80'h001084ce994fab5e6ffe;
mem[6890] = 80'h0110ce437f4c40581cfa;
mem[6891] = 80'h00000000000000000000;
mem[6892] = 80'h10100000010000010010;
mem[6893] = 80'h00109400000208004500;
mem[6894] = 80'h0010002e2b710000fffd;
mem[6895] = 80'h00100e09c0550102c000;
mem[6896] = 80'h00100001ffabffabffab;
mem[6897] = 80'h00108ef167c3cef0da44;
mem[6898] = 80'h00104f1c1ea25e8e2eaf;
mem[6899] = 80'h01108174e3a4ffb3f20a;
mem[6900] = 80'h00000000000000000000;
mem[6901] = 80'h00000000000000000000;
mem[6902] = 80'h00000000000000000000;
mem[6903] = 80'h00000000000000000000;
mem[6904] = 80'h10100000010000010010;
mem[6905] = 80'h00109400000208004500;
mem[6906] = 80'h0010002e2b720000fffd;
mem[6907] = 80'h00100e08c0550102c000;
mem[6908] = 80'h00100001ffabffabffab;
mem[6909] = 80'h00108d6305b6a67a9d84;
mem[6910] = 80'h0010136b969440fe9d5d;
mem[6911] = 80'h011048555836f475bf1a;
mem[6912] = 80'h00000000000000000000;
mem[6913] = 80'h10100000010000010010;
mem[6914] = 80'h00109400000208004500;
mem[6915] = 80'h0010002e2b730000fffd;
mem[6916] = 80'h00100e07c0550102c000;
mem[6917] = 80'h00100001ffabffabffab;
mem[6918] = 80'h00108c12db9a7e035f3b;
mem[6919] = 80'h0010d8b91179b52e9e0c;
mem[6920] = 80'h01106ccc10d95b52efae;
mem[6921] = 80'h00000000000000000000;
mem[6922] = 80'h00000000000000000000;
mem[6923] = 80'h00000000000000000000;
mem[6924] = 80'h00000000000000000000;
mem[6925] = 80'h10100000010000010010;
mem[6926] = 80'h00109400000208004500;
mem[6927] = 80'h0010002e2b740000fffd;
mem[6928] = 80'h00100e06c0550102c000;
mem[6929] = 80'h00100001ffabffabffab;
mem[6930] = 80'h00108b361f70af17d0bb;
mem[6931] = 80'h00106056001589cfede9;
mem[6932] = 80'h0110749988c732c116cd;
mem[6933] = 80'h00000000000000000000;
mem[6934] = 80'h00000000000000000000;
mem[6935] = 80'h00000000000000000000;
mem[6936] = 80'h10100000010000010010;
mem[6937] = 80'h00109400000208004500;
mem[6938] = 80'h0010002e2b750000fffd;
mem[6939] = 80'h00100e05c0550102c000;
mem[6940] = 80'h00100001ffabffabffab;
mem[6941] = 80'h00108a47c15c776e1204;
mem[6942] = 80'h0010ab8487f87c1e72b8;
mem[6943] = 80'h01103ab6cdde17757283;
mem[6944] = 80'h00000000000000000000;
mem[6945] = 80'h10100000010000010010;
mem[6946] = 80'h00109400000208004500;
mem[6947] = 80'h0010002e2b760000fffd;
mem[6948] = 80'h00100e04c0550102c000;
mem[6949] = 80'h00100001ffabffabffab;
mem[6950] = 80'h001089d5a3291fe455c4;
mem[6951] = 80'h0010f7f30fce626ef94a;
mem[6952] = 80'h01107fab7a312661e973;
mem[6953] = 80'h00000000000000000000;
mem[6954] = 80'h00000000000000000000;
mem[6955] = 80'h00000000000000000000;
mem[6956] = 80'h00000000000000000000;
mem[6957] = 80'h10100000010000010010;
mem[6958] = 80'h00109400000208004500;
mem[6959] = 80'h0010002e2b770000fffd;
mem[6960] = 80'h00100e03c0550102c000;
mem[6961] = 80'h00100001ffabffabffab;
mem[6962] = 80'h001088a47d05c79d977b;
mem[6963] = 80'h00103c21882397bef21b;
mem[6964] = 80'h0110d29b7a81d7732364;
mem[6965] = 80'h00000000000000000000;
mem[6966] = 80'h00000000000000000000;
mem[6967] = 80'h00000000000000000000;
mem[6968] = 80'h10100000010000010010;
mem[6969] = 80'h00109400000208004500;
mem[6970] = 80'h0010002e2b780000fffd;
mem[6971] = 80'h00100e02c0550102c000;
mem[6972] = 80'h00100001ffabffabffab;
mem[6973] = 80'h0010879c2afcbdcd4ac5;
mem[6974] = 80'h0010862d2d161bac0d81;
mem[6975] = 80'h011009005f63832f2a80;
mem[6976] = 80'h00000000000000000000;
mem[6977] = 80'h10100000010000010010;
mem[6978] = 80'h00109400000208004500;
mem[6979] = 80'h0010002e2b790000fffd;
mem[6980] = 80'h00100e01c0550102c000;
mem[6981] = 80'h00100001ffabffabffab;
mem[6982] = 80'h001086edf4d065b4887a;
mem[6983] = 80'h00104dffaafbee7c73d0;
mem[6984] = 80'h0110539ce72d13835ff9;
mem[6985] = 80'h00000000000000000000;
mem[6986] = 80'h00000000000000000000;
mem[6987] = 80'h00000000000000000000;
mem[6988] = 80'h10100000010000010010;
mem[6989] = 80'h00109400000208004500;
mem[6990] = 80'h0010002e2b7a0000fffd;
mem[6991] = 80'h00100e00c0550102c000;
mem[6992] = 80'h00100001ffabffabffab;
mem[6993] = 80'h0010857f96a50d3ecfba;
mem[6994] = 80'h0010118822cdf00c3122;
mem[6995] = 80'h0110ba4df70fe485b8a4;
mem[6996] = 80'h00000000000000000000;
mem[6997] = 80'h00000000000000000000;
mem[6998] = 80'h00000000000000000000;
mem[6999] = 80'h10100000010000010010;
mem[7000] = 80'h00109400000208004500;
mem[7001] = 80'h0010002e2b7b0000fffd;
mem[7002] = 80'h00100dffc0550102c000;
mem[7003] = 80'h00100001ffabffabffab;
mem[7004] = 80'h0010840e4889d5470d05;
mem[7005] = 80'h0010da5aa52005dc7273;
mem[7006] = 80'h01109318c637c31212d1;
mem[7007] = 80'h00000000000000000000;
mem[7008] = 80'h10100000010000010010;
mem[7009] = 80'h00109400000208004500;
mem[7010] = 80'h0010002e2b7c0000fffd;
mem[7011] = 80'h00100dfec0550102c000;
mem[7012] = 80'h00100001ffabffabffab;
mem[7013] = 80'h0010832a8c6304538285;
mem[7014] = 80'h001062b5b44c393d5196;
mem[7015] = 80'h011085f241d1f33384ee;
mem[7016] = 80'h00000000000000000000;
mem[7017] = 80'h00000000000000000000;
mem[7018] = 80'h00000000000000000000;
mem[7019] = 80'h00000000000000000000;
mem[7020] = 80'h10100000010000010010;
mem[7021] = 80'h00109400000208004500;
mem[7022] = 80'h0010002e2b7d0000fffd;
mem[7023] = 80'h00100dfdc0550102c000;
mem[7024] = 80'h00100001ffabffabffab;
mem[7025] = 80'h0010825b524fdc2a403a;
mem[7026] = 80'h0010a96733a1cced1ec7;
mem[7027] = 80'h0110e9ca5c67282bf033;
mem[7028] = 80'h00000000000000000000;
mem[7029] = 80'h00000000000000000000;
mem[7030] = 80'h00000000000000000000;
mem[7031] = 80'h10100000010000010010;
mem[7032] = 80'h00109400000208004500;
mem[7033] = 80'h0010002e2b7e0000fffd;
mem[7034] = 80'h00100dfcc0550102c000;
mem[7035] = 80'h00100001ffabffabffab;
mem[7036] = 80'h001081c9303ab4a007fa;
mem[7037] = 80'h0010f510bb97d29e5535;
mem[7038] = 80'h0110e3d3d5108cdb0498;
mem[7039] = 80'h00000000000000000000;
mem[7040] = 80'h10100000010000010010;
mem[7041] = 80'h00109400000208004500;
mem[7042] = 80'h0010002e2b7f0000fffd;
mem[7043] = 80'h00100dfbc0550102c000;
mem[7044] = 80'h00100001ffabffabffab;
mem[7045] = 80'h001080b8ee166cd9c545;
mem[7046] = 80'h00103ec23c7a274e2c64;
mem[7047] = 80'h011020d86f4aa2a21664;
mem[7048] = 80'h00000000000000000000;
mem[7049] = 80'h00000000000000000000;
mem[7050] = 80'h00000000000000000000;
mem[7051] = 80'h00000000000000000000;
mem[7052] = 80'h10100000010000010010;
mem[7053] = 80'h00109400000208004500;
mem[7054] = 80'h0010002e2b800000fffd;
mem[7055] = 80'h00100dfac0550102c000;
mem[7056] = 80'h00100001ffabffabffab;
mem[7057] = 80'h00107f97a40ddb0e84d0;
mem[7058] = 80'h0010787341217401d6ab;
mem[7059] = 80'h011097eae04e57bb5be7;
mem[7060] = 80'h00000000000000000000;
mem[7061] = 80'h10100000010000010010;
mem[7062] = 80'h00109400000208004500;
mem[7063] = 80'h0010002e2b810000fffd;
mem[7064] = 80'h00100df9c0550102c000;
mem[7065] = 80'h00100001ffabffabffab;
mem[7066] = 80'h00107ee67a210377466f;
mem[7067] = 80'h0010b3a1c6cc81d1dffa;
mem[7068] = 80'h01105cb8841e45a046c1;
mem[7069] = 80'h00000000000000000000;
mem[7070] = 80'h00000000000000000000;
mem[7071] = 80'h00000000000000000000;
mem[7072] = 80'h00000000000000000000;
mem[7073] = 80'h10100000010000010010;
mem[7074] = 80'h00109400000208004500;
mem[7075] = 80'h0010002e2b820000fffd;
mem[7076] = 80'h00100df8c0550102c000;
mem[7077] = 80'h00100001ffabffabffab;
mem[7078] = 80'h00107d7418546bfd01af;
mem[7079] = 80'h0010efd64efa9fa14a08;
mem[7080] = 80'h011039d99a3626b91d8f;
mem[7081] = 80'h00000000000000000000;
mem[7082] = 80'h00000000000000000000;
mem[7083] = 80'h00000000000000000000;
mem[7084] = 80'h10100000010000010010;
mem[7085] = 80'h00109400000208004500;
mem[7086] = 80'h0010002e2b830000fffd;
mem[7087] = 80'h00100df7c0550102c000;
mem[7088] = 80'h00100001ffabffabffab;
mem[7089] = 80'h00107c05c678b384c310;
mem[7090] = 80'h00102404c9176a71c859;
mem[7091] = 80'h011035e9f11b376c4d96;
mem[7092] = 80'h00000000000000000000;
mem[7093] = 80'h10100000010000010010;
mem[7094] = 80'h00109400000208004500;
mem[7095] = 80'h0010002e2b840000fffd;
mem[7096] = 80'h00100df6c0550102c000;
mem[7097] = 80'h00100001ffabffabffab;
mem[7098] = 80'h00107b21029262904c90;
mem[7099] = 80'h00109cebd87b5690babc;
mem[7100] = 80'h01101e8d2deafb817f5d;
mem[7101] = 80'h00000000000000000000;
mem[7102] = 80'h00000000000000000000;
mem[7103] = 80'h00000000000000000000;
mem[7104] = 80'h00000000000000000000;
mem[7105] = 80'h10100000010000010010;
mem[7106] = 80'h00109400000208004500;
mem[7107] = 80'h0010002e2b850000fffd;
mem[7108] = 80'h00100df5c0550102c000;
mem[7109] = 80'h00100001ffabffabffab;
mem[7110] = 80'h00107a50dcbebae98e2f;
mem[7111] = 80'h001057395f96a340c4ed;
mem[7112] = 80'h01104411fcc767cd8e44;
mem[7113] = 80'h00000000000000000000;
mem[7114] = 80'h10100000010000010010;
mem[7115] = 80'h00109400000208004500;
mem[7116] = 80'h0010002e2b860000fffd;
mem[7117] = 80'h00100df4c0550102c000;
mem[7118] = 80'h00100001ffabffabffab;
mem[7119] = 80'h001079c2becbd263c9ef;
mem[7120] = 80'h00100b4ed7a0bd300d1f;
mem[7121] = 80'h01106aa2133dee41fbd6;
mem[7122] = 80'h00000000000000000000;
mem[7123] = 80'h00000000000000000000;
mem[7124] = 80'h00000000000000000000;
mem[7125] = 80'h00000000000000000000;
mem[7126] = 80'h10100000010000010010;
mem[7127] = 80'h00109400000208004500;
mem[7128] = 80'h0010002e2b870000fffd;
mem[7129] = 80'h00100df3c0550102c000;
mem[7130] = 80'h00100001ffabffabffab;
mem[7131] = 80'h001078b360e70a1a0b50;
mem[7132] = 80'h0010c09c504d48e0444e;
mem[7133] = 80'h0110ac3cc6a5b0619a75;
mem[7134] = 80'h00000000000000000000;
mem[7135] = 80'h00000000000000000000;
mem[7136] = 80'h00000000000000000000;
mem[7137] = 80'h10100000010000010010;
mem[7138] = 80'h00109400000208004500;
mem[7139] = 80'h0010002e2b880000fffd;
mem[7140] = 80'h00100df2c0550102c000;
mem[7141] = 80'h00100001ffabffabffab;
mem[7142] = 80'h0010778b371e704ad6ee;
mem[7143] = 80'h00107a90f578c4f364d4;
mem[7144] = 80'h0110458e2abdeaa262fe;
mem[7145] = 80'h00000000000000000000;
mem[7146] = 80'h10100000010000010010;
mem[7147] = 80'h00109400000208004500;
mem[7148] = 80'h0010002e2b890000fffd;
mem[7149] = 80'h00100df1c0550102c000;
mem[7150] = 80'h00100001ffabffabffab;
mem[7151] = 80'h001076fae932a8331451;
mem[7152] = 80'h0010b142729531232585;
mem[7153] = 80'h01100ab95e14b741f099;
mem[7154] = 80'h00000000000000000000;
mem[7155] = 80'h00000000000000000000;
mem[7156] = 80'h00000000000000000000;
mem[7157] = 80'h00000000000000000000;
mem[7158] = 80'h10100000010000010010;
mem[7159] = 80'h00109400000208004500;
mem[7160] = 80'h0010002e2b8a0000fffd;
mem[7161] = 80'h00100df0c0550102c000;
mem[7162] = 80'h00100001ffabffabffab;
mem[7163] = 80'h001075688b47c0b95391;
mem[7164] = 80'h0010ed35faa32f53e677;
mem[7165] = 80'h0110cbc1219eb13dbc98;
mem[7166] = 80'h00000000000000000000;
mem[7167] = 80'h10100000010000010010;
mem[7168] = 80'h00109400000208004500;
mem[7169] = 80'h0010002e2b8b0000fffd;
mem[7170] = 80'h00100defc0550102c000;
mem[7171] = 80'h00100001ffabffabffab;
mem[7172] = 80'h00107419556b18c0912e;
mem[7173] = 80'h001026e77d4eda83a526;
mem[7174] = 80'h0110e29486178ec8a67b;
mem[7175] = 80'h00000000000000000000;
mem[7176] = 80'h00000000000000000000;
mem[7177] = 80'h00000000000000000000;
mem[7178] = 80'h00000000000000000000;
mem[7179] = 80'h10100000010000010010;
mem[7180] = 80'h00109400000208004500;
mem[7181] = 80'h0010002e2b8c0000fffd;
mem[7182] = 80'h00100deec0550102c000;
mem[7183] = 80'h00100001ffabffabffab;
mem[7184] = 80'h0010733d9181c9d41eae;
mem[7185] = 80'h00109e086c22e662e7c3;
mem[7186] = 80'h0110cc656e0649b9c863;
mem[7187] = 80'h00000000000000000000;
mem[7188] = 80'h00000000000000000000;
mem[7189] = 80'h00000000000000000000;
mem[7190] = 80'h10100000010000010010;
mem[7191] = 80'h00109400000208004500;
mem[7192] = 80'h0010002e2b8d0000fffd;
mem[7193] = 80'h00100dedc0550102c000;
mem[7194] = 80'h00100001ffabffabffab;
mem[7195] = 80'h0010724c4fad11addc11;
mem[7196] = 80'h001055daebcf13b26992;
mem[7197] = 80'h011085380c2039cc50e5;
mem[7198] = 80'h00000000000000000000;
mem[7199] = 80'h10100000010000010010;
mem[7200] = 80'h00109400000208004500;
mem[7201] = 80'h0010002e2b8e0000fffd;
mem[7202] = 80'h00100decc0550102c000;
mem[7203] = 80'h00100001ffabffabffab;
mem[7204] = 80'h001071de2dd879279bd1;
mem[7205] = 80'h001009ad63f90dc2e360;
mem[7206] = 80'h0110f314f971496036f7;
mem[7207] = 80'h00000000000000000000;
mem[7208] = 80'h00000000000000000000;
mem[7209] = 80'h00000000000000000000;
mem[7210] = 80'h10100000010000010010;
mem[7211] = 80'h00109400000208004500;
mem[7212] = 80'h0010002e2b8f0000fffd;
mem[7213] = 80'h00100debc0550102c000;
mem[7214] = 80'h00100001ffabffabffab;
mem[7215] = 80'h001070aff3f4a15e596e;
mem[7216] = 80'h0010c27fe414f812f831;
mem[7217] = 80'h01105d57ac5dba7f5d99;
mem[7218] = 80'h00000000000000000000;
mem[7219] = 80'h00000000000000000000;
mem[7220] = 80'h00000000000000000000;
mem[7221] = 80'h10100000010000010010;
mem[7222] = 80'h00109400000208004500;
mem[7223] = 80'h0010002e2b900000fffd;
mem[7224] = 80'h00100deac0550102c000;
mem[7225] = 80'h00100001ffabffabffab;
mem[7226] = 80'h00106fae822a8d8620ac;
mem[7227] = 80'h00107db4299215e70c54;
mem[7228] = 80'h011057703f02bd8c3090;
mem[7229] = 80'h00000000000000000000;
mem[7230] = 80'h00000000000000000000;
mem[7231] = 80'h00000000000000000000;
mem[7232] = 80'h10100000010000010010;
mem[7233] = 80'h00109400000208004500;
mem[7234] = 80'h0010002e2b910000fffd;
mem[7235] = 80'h00100de9c0550102c000;
mem[7236] = 80'h00100001ffabffabffab;
mem[7237] = 80'h00106edf5c0655ffe213;
mem[7238] = 80'h0010b666ae7fe0388305;
mem[7239] = 80'h0110012d33b5b3f8b05f;
mem[7240] = 80'h00000000000000000000;
mem[7241] = 80'h10100000010000010010;
mem[7242] = 80'h00109400000208004500;
mem[7243] = 80'h0010002e2b920000fffd;
mem[7244] = 80'h00100de8c0550102c000;
mem[7245] = 80'h00100001ffabffabffab;
mem[7246] = 80'h00106d4d3e733d75a5d3;
mem[7247] = 80'h0010ea112649fe4830f7;
mem[7248] = 80'h0110c80c694ee925f63c;
mem[7249] = 80'h00000000000000000000;
mem[7250] = 80'h00000000000000000000;
mem[7251] = 80'h00000000000000000000;
mem[7252] = 80'h10100000010000010010;
mem[7253] = 80'h00109400000208004500;
mem[7254] = 80'h0010002e2b930000fffd;
mem[7255] = 80'h00100de7c0550102c000;
mem[7256] = 80'h00100001ffabffabffab;
mem[7257] = 80'h00106c3ce05fe50c676c;
mem[7258] = 80'h001021c3a1a40b9873a6;
mem[7259] = 80'h0110e15942eaaf1fff42;
mem[7260] = 80'h00000000000000000000;
mem[7261] = 80'h00000000000000000000;
mem[7262] = 80'h00000000000000000000;
mem[7263] = 80'h10100000010000010010;
mem[7264] = 80'h00109400000208004500;
mem[7265] = 80'h0010002e2b940000fffd;
mem[7266] = 80'h00100de6c0550102c000;
mem[7267] = 80'h00100001ffabffabffab;
mem[7268] = 80'h00106b1824b53418e8ec;
mem[7269] = 80'h0010992cb0c837794043;
mem[7270] = 80'h0110f4c09cba47b5c673;
mem[7271] = 80'h00000000000000000000;
mem[7272] = 80'h00000000000000000000;
mem[7273] = 80'h00000000000000000000;
mem[7274] = 80'h10100000010000010010;
mem[7275] = 80'h00109400000208004500;
mem[7276] = 80'h0010002e2b950000fffd;
mem[7277] = 80'h00100de5c0550102c000;
mem[7278] = 80'h00100001ffabffabffab;
mem[7279] = 80'h00106a69fa99ec612a53;
mem[7280] = 80'h001052fe3725c2a90112;
mem[7281] = 80'h0110bbf77a70608e9883;
mem[7282] = 80'h00000000000000000000;
mem[7283] = 80'h10100000010000010010;
mem[7284] = 80'h00109400000208004500;
mem[7285] = 80'h0010002e2b960000fffd;
mem[7286] = 80'h00100de4c0550102c000;
mem[7287] = 80'h00100001ffabffabffab;
mem[7288] = 80'h001069fb98ec84eb6d93;
mem[7289] = 80'h00100e89bf13dcd954e0;
mem[7290] = 80'h0110c8c2427fd73138a4;
mem[7291] = 80'h00000000000000000000;
mem[7292] = 80'h00000000000000000000;
mem[7293] = 80'h00000000000000000000;
mem[7294] = 80'h00000000000000000000;
mem[7295] = 80'h10100000010000010010;
mem[7296] = 80'h00109400000208004500;
mem[7297] = 80'h0010002e2b970000fffd;
mem[7298] = 80'h00100de3c0550102c000;
mem[7299] = 80'h00100001ffabffabffab;
mem[7300] = 80'h0010688a46c05c92af2c;
mem[7301] = 80'h0010c55b38fe29091eb1;
mem[7302] = 80'h01105b0fa3d28a3b7dfe;
mem[7303] = 80'h00000000000000000000;
mem[7304] = 80'h00000000000000000000;
mem[7305] = 80'h00000000000000000000;
mem[7306] = 80'h10100000010000010010;
mem[7307] = 80'h00109400000208004500;
mem[7308] = 80'h0010002e2b980000fffd;
mem[7309] = 80'h00100de2c0550102c000;
mem[7310] = 80'h00100001ffabffabffab;
mem[7311] = 80'h001067b2113926c27292;
mem[7312] = 80'h00107f579dcba51ba12b;
mem[7313] = 80'h01108d58fcfcacc5f138;
mem[7314] = 80'h00000000000000000000;
mem[7315] = 80'h10100000010000010010;
mem[7316] = 80'h00109400000208004500;
mem[7317] = 80'h0010002e2b990000fffd;
mem[7318] = 80'h00100de1c0550102c000;
mem[7319] = 80'h00100001ffabffabffab;
mem[7320] = 80'h001066c3cf15febbb02d;
mem[7321] = 80'h0010b4851a2650cbdf7a;
mem[7322] = 80'h0110d7c44486899d3060;
mem[7323] = 80'h00000000000000000000;
mem[7324] = 80'h00000000000000000000;
mem[7325] = 80'h00000000000000000000;
mem[7326] = 80'h10100000010000010010;
mem[7327] = 80'h00109400000208004500;
mem[7328] = 80'h0010002e2b9a0000fffd;
mem[7329] = 80'h00100de0c0550102c000;
mem[7330] = 80'h00100001ffabffabffab;
mem[7331] = 80'h00106551ad609631f7ed;
mem[7332] = 80'h0010e8f292104ebb5e88;
mem[7333] = 80'h01107d12b9d4afea909d;
mem[7334] = 80'h00000000000000000000;
mem[7335] = 80'h00000000000000000000;
mem[7336] = 80'h00000000000000000000;
mem[7337] = 80'h10100000010000010010;
mem[7338] = 80'h00109400000208004500;
mem[7339] = 80'h0010002e2b9b0000fffd;
mem[7340] = 80'h00100ddfc0550102c000;
mem[7341] = 80'h00100001ffabffabffab;
mem[7342] = 80'h00106420734c4e483552;
mem[7343] = 80'h0010232015fdbb6adfd9;
mem[7344] = 80'h01101341bd5523589692;
mem[7345] = 80'h00000000000000000000;
mem[7346] = 80'h00000000000000000000;
mem[7347] = 80'h00000000000000000000;
mem[7348] = 80'h10100000010000010010;
mem[7349] = 80'h00109400000208004500;
mem[7350] = 80'h0010002e2b9c0000fffd;
mem[7351] = 80'h00100ddec0550102c000;
mem[7352] = 80'h00100001ffabffabffab;
mem[7353] = 80'h00106304b7a69f5cbad2;
mem[7354] = 80'h00109bcf0491878bba3c;
mem[7355] = 80'h0110a2c1063bc58d6d71;
mem[7356] = 80'h00000000000000000000;
mem[7357] = 80'h10100000010000010010;
mem[7358] = 80'h00109400000208004500;
mem[7359] = 80'h0010002e2b9d0000fffd;
mem[7360] = 80'h00100dddc0550102c000;
mem[7361] = 80'h00100001ffabffabffab;
mem[7362] = 80'h00106275698a4725786d;
mem[7363] = 80'h0010501d837c725bb36d;
mem[7364] = 80'h011069931177ade06347;
mem[7365] = 80'h00000000000000000000;
mem[7366] = 80'h00000000000000000000;
mem[7367] = 80'h00000000000000000000;
mem[7368] = 80'h10100000010000010010;
mem[7369] = 80'h00109400000208004500;
mem[7370] = 80'h0010002e2b9e0000fffd;
mem[7371] = 80'h00100ddcc0550102c000;
mem[7372] = 80'h00100001ffabffabffab;
mem[7373] = 80'h001061e70bff2faf3fad;
mem[7374] = 80'h00100c6a0b4a6c2b3a9f;
mem[7375] = 80'h01104aec1952df7bc2b7;
mem[7376] = 80'h00000000000000000000;
mem[7377] = 80'h00000000000000000000;
mem[7378] = 80'h00000000000000000000;
mem[7379] = 80'h10100000010000010010;
mem[7380] = 80'h00109400000208004500;
mem[7381] = 80'h0010002e2b9f0000fffd;
mem[7382] = 80'h00100ddbc0550102c000;
mem[7383] = 80'h00100001ffabffabffab;
mem[7384] = 80'h00106096d5d3f7d6fd12;
mem[7385] = 80'h0010c7b88ca799fb42ce;
mem[7386] = 80'h0110bad6e8aab65dee6c;
mem[7387] = 80'h00000000000000000000;
mem[7388] = 80'h00000000000000000000;
mem[7389] = 80'h00000000000000000000;
mem[7390] = 80'h10100000010000010010;
mem[7391] = 80'h00109400000208004500;
mem[7392] = 80'h0010002e2ba00000fffd;
mem[7393] = 80'h00100ddac0550102c000;
mem[7394] = 80'h00100001ffabffabffab;
mem[7395] = 80'h00105fe5e843761fcc28;
mem[7396] = 80'h001073fd9047b7c06c55;
mem[7397] = 80'h011063a0e99221d3a6df;
mem[7398] = 80'h00000000000000000000;
mem[7399] = 80'h10100000010000010010;
mem[7400] = 80'h00109400000208004500;
mem[7401] = 80'h0010002e2ba10000fffd;
mem[7402] = 80'h00100dd9c0550102c000;
mem[7403] = 80'h00100001ffabffabffab;
mem[7404] = 80'h00105e94366fae660e97;
mem[7405] = 80'h0010b82f17aa42102d04;
mem[7406] = 80'h01102c97427910c94626;
mem[7407] = 80'h00000000000000000000;
mem[7408] = 80'h00000000000000000000;
mem[7409] = 80'h00000000000000000000;
mem[7410] = 80'h00000000000000000000;
mem[7411] = 80'h10100000010000010010;
mem[7412] = 80'h00109400000208004500;
mem[7413] = 80'h0010002e2ba20000fffd;
mem[7414] = 80'h00100dd8c0550102c000;
mem[7415] = 80'h00100001ffabffabffab;
mem[7416] = 80'h00105d06541ac6ec4957;
mem[7417] = 80'h0010e4589f9c5c60fff6;
mem[7418] = 80'h0110ddad80a09c15bccf;
mem[7419] = 80'h00000000000000000000;
mem[7420] = 80'h00000000000000000000;
mem[7421] = 80'h00000000000000000000;
mem[7422] = 80'h10100000010000010010;
mem[7423] = 80'h00109400000208004500;
mem[7424] = 80'h0010002e2ba30000fffd;
mem[7425] = 80'h00100dd7c0550102c000;
mem[7426] = 80'h00100001ffabffabffab;
mem[7427] = 80'h00105c778a361e958be8;
mem[7428] = 80'h00102f8a1871a9b0bda7;
mem[7429] = 80'h0110c7c9f7b66fe4bf8e;
mem[7430] = 80'h00000000000000000000;
mem[7431] = 80'h10100000010000010010;
mem[7432] = 80'h00109400000208004500;
mem[7433] = 80'h0010002e2ba40000fffd;
mem[7434] = 80'h00100dd6c0550102c000;
mem[7435] = 80'h00100001ffabffabffab;
mem[7436] = 80'h00105b534edccf810468;
mem[7437] = 80'h00109765091d95520f42;
mem[7438] = 80'h0110a3a999257321bcd4;
mem[7439] = 80'h00000000000000000000;
mem[7440] = 80'h00000000000000000000;
mem[7441] = 80'h00000000000000000000;
mem[7442] = 80'h10100000010000010010;
mem[7443] = 80'h00109400000208004500;
mem[7444] = 80'h0010002e2ba50000fffd;
mem[7445] = 80'h00100dd5c0550102c000;
mem[7446] = 80'h00100001ffabffabffab;
mem[7447] = 80'h00105a2290f017f8c6d7;
mem[7448] = 80'h00105cb78ef060827013;
mem[7449] = 80'h0110ca04afda71b0c4b8;
mem[7450] = 80'h00000000000000000000;
mem[7451] = 80'h00000000000000000000;
mem[7452] = 80'h00000000000000000000;
mem[7453] = 80'h10100000010000010010;
mem[7454] = 80'h00109400000208004500;
mem[7455] = 80'h0010002e2ba60000fffd;
mem[7456] = 80'h00100dd4c0550102c000;
mem[7457] = 80'h00100001ffabffabffab;
mem[7458] = 80'h001059b0f2857f728117;
mem[7459] = 80'h001000c006c67ef2fbe1;
mem[7460] = 80'h01108f19a1cbaa6e5d27;
mem[7461] = 80'h00000000000000000000;
mem[7462] = 80'h00000000000000000000;
mem[7463] = 80'h00000000000000000000;
mem[7464] = 80'h10100000010000010010;
mem[7465] = 80'h00109400000208004500;
mem[7466] = 80'h0010002e2ba70000fffd;
mem[7467] = 80'h00100dd3c0550102c000;
mem[7468] = 80'h00100001ffabffabffab;
mem[7469] = 80'h001058c12ca9a70b43a8;
mem[7470] = 80'h0010cb12812b8b22f0b0;
mem[7471] = 80'h01102229a5a6361799ac;
mem[7472] = 80'h00000000000000000000;
mem[7473] = 80'h10100000010000010010;
mem[7474] = 80'h00109400000208004500;
mem[7475] = 80'h0010002e2ba80000fffd;
mem[7476] = 80'h00100dd2c0550102c000;
mem[7477] = 80'h00100001ffabffabffab;
mem[7478] = 80'h001057f97b50dd5b9e16;
mem[7479] = 80'h0010711e241e07300e2a;
mem[7480] = 80'h0110ca833c297ebc883f;
mem[7481] = 80'h00000000000000000000;
mem[7482] = 80'h00000000000000000000;
mem[7483] = 80'h00000000000000000000;
mem[7484] = 80'h10100000010000010010;
mem[7485] = 80'h00109400000208004500;
mem[7486] = 80'h0010002e2ba90000fffd;
mem[7487] = 80'h00100dd1c0550102c000;
mem[7488] = 80'h00100001ffabffabffab;
mem[7489] = 80'h00105688a57c05225ca9;
mem[7490] = 80'h0010bacca3f3f2e0917b;
mem[7491] = 80'h0110b39c0b76b6d9ba1c;
mem[7492] = 80'h00000000000000000000;
mem[7493] = 80'h00000000000000000000;
mem[7494] = 80'h00000000000000000000;
mem[7495] = 80'h10100000010000010010;
mem[7496] = 80'h00109400000208004500;
mem[7497] = 80'h0010002e2baa0000fffd;
mem[7498] = 80'h00100dd0c0550102c000;
mem[7499] = 80'h00100001ffabffabffab;
mem[7500] = 80'h0010551ac7096da81b69;
mem[7501] = 80'h0010e6bb2bc5ec901189;
mem[7502] = 80'h01102a7b1fb43c7ec292;
mem[7503] = 80'h00000000000000000000;
mem[7504] = 80'h00000000000000000000;
mem[7505] = 80'h00000000000000000000;
mem[7506] = 80'h10100000010000010010;
mem[7507] = 80'h00109400000208004500;
mem[7508] = 80'h0010002e2bab0000fffd;
mem[7509] = 80'h00100dcfc0550102c000;
mem[7510] = 80'h00100001ffabffabffab;
mem[7511] = 80'h0010546b1925b5d1d9d6;
mem[7512] = 80'h00102d69ac28194011d8;
mem[7513] = 80'h01105bb1a26b5b25c732;
mem[7514] = 80'h00000000000000000000;
mem[7515] = 80'h10100000010000010010;
mem[7516] = 80'h00109400000208004500;
mem[7517] = 80'h0010002e2bac0000fffd;
mem[7518] = 80'h00100dcec0550102c000;
mem[7519] = 80'h00100001ffabffabffab;
mem[7520] = 80'h0010534fddcf64c55656;
mem[7521] = 80'h00109586bd4425a1553d;
mem[7522] = 80'h0110dfe666340b6886ab;
mem[7523] = 80'h00000000000000000000;
mem[7524] = 80'h00000000000000000000;
mem[7525] = 80'h00000000000000000000;
mem[7526] = 80'h00000000000000000000;
mem[7527] = 80'h10100000010000010010;
mem[7528] = 80'h00109400000208004500;
mem[7529] = 80'h0010002e2bad0000fffd;
mem[7530] = 80'h00100dcdc0550102c000;
mem[7531] = 80'h00100001ffabffabffab;
mem[7532] = 80'h0010523e03e3bcbc94e9;
mem[7533] = 80'h00105e543aa9d0711c6c;
mem[7534] = 80'h01101978b8e49e0b8e1b;
mem[7535] = 80'h00000000000000000000;
mem[7536] = 80'h00000000000000000000;
mem[7537] = 80'h00000000000000000000;
mem[7538] = 80'h10100000010000010010;
mem[7539] = 80'h00109400000208004500;
mem[7540] = 80'h0010002e2bae0000fffd;
mem[7541] = 80'h00100dccc0550102c000;
mem[7542] = 80'h00100001ffabffabffab;
mem[7543] = 80'h001051ac6196d436d329;
mem[7544] = 80'h00100223b29fce00569e;
mem[7545] = 80'h01104e307dca1743dbf6;
mem[7546] = 80'h00000000000000000000;
mem[7547] = 80'h10100000010000010010;
mem[7548] = 80'h00109400000208004500;
mem[7549] = 80'h0010002e2baf0000fffd;
mem[7550] = 80'h00100dcbc0550102c000;
mem[7551] = 80'h00100001ffabffabffab;
mem[7552] = 80'h001050ddbfba0c4f1196;
mem[7553] = 80'h0010c9f135723bd00ccf;
mem[7554] = 80'h0110de8eaaf0a4a53d0c;
mem[7555] = 80'h00000000000000000000;
mem[7556] = 80'h00000000000000000000;
mem[7557] = 80'h00000000000000000000;
mem[7558] = 80'h10100000010000010010;
mem[7559] = 80'h00109400000208004500;
mem[7560] = 80'h0010002e2bb00000fffd;
mem[7561] = 80'h00100dcac0550102c000;
mem[7562] = 80'h00100001ffabffabffab;
mem[7563] = 80'h00104fdcce6420976854;
mem[7564] = 80'h0010763af8f4d625b6aa;
mem[7565] = 80'h0110fa6a6268271e49bf;
mem[7566] = 80'h00000000000000000000;
mem[7567] = 80'h10100000010000010010;
mem[7568] = 80'h00109400000208004500;
mem[7569] = 80'h0010002e2bb10000fffd;
mem[7570] = 80'h00100dc9c0550102c000;
mem[7571] = 80'h00100001ffabffabffab;
mem[7572] = 80'h00104ead1048f8eeaaeb;
mem[7573] = 80'h0010bde87f1923f5f7fb;
mem[7574] = 80'h0110b55deede3a9bb689;
mem[7575] = 80'h00000000000000000000;
mem[7576] = 80'h00000000000000000000;
mem[7577] = 80'h00000000000000000000;
mem[7578] = 80'h00000000000000000000;
mem[7579] = 80'h10100000010000010010;
mem[7580] = 80'h00109400000208004500;
mem[7581] = 80'h0010002e2bb20000fffd;
mem[7582] = 80'h00100dc8c0550102c000;
mem[7583] = 80'h00100001ffabffabffab;
mem[7584] = 80'h00104d3f723d9064ed2b;
mem[7585] = 80'h0010e19ff72f3d854609;
mem[7586] = 80'h01101a1e4c76013b21dc;
mem[7587] = 80'h00000000000000000000;
mem[7588] = 80'h00000000000000000000;
mem[7589] = 80'h00000000000000000000;
mem[7590] = 80'h10100000010000010010;
mem[7591] = 80'h00109400000208004500;
mem[7592] = 80'h0010002e2bb30000fffd;
mem[7593] = 80'h00100dc7c0550102c000;
mem[7594] = 80'h00100001ffabffabffab;
mem[7595] = 80'h00104c4eac11481d2f94;
mem[7596] = 80'h00102a4d70c2c855c758;
mem[7597] = 80'h0110437d21b30b3e4729;
mem[7598] = 80'h00000000000000000000;
mem[7599] = 80'h00000000000000000000;
mem[7600] = 80'h00000000000000000000;
mem[7601] = 80'h10100000010000010010;
mem[7602] = 80'h00109400000208004500;
mem[7603] = 80'h0010002e2bb40000fffd;
mem[7604] = 80'h00100dc6c0550102c000;
mem[7605] = 80'h00100001ffabffabffab;
mem[7606] = 80'h00104b6a68fb9909a014;
mem[7607] = 80'h001092a261aef4b4b2bd;
mem[7608] = 80'h0110f18e85290aa8e2fa;
mem[7609] = 80'h00000000000000000000;
mem[7610] = 80'h10100000010000010010;
mem[7611] = 80'h00109400000208004500;
mem[7612] = 80'h0010002e2bb50000fffd;
mem[7613] = 80'h00100dc5c0550102c000;
mem[7614] = 80'h00100001ffabffabffab;
mem[7615] = 80'h00104a1bb6d7417062ab;
mem[7616] = 80'h00105970e6430164aaec;
mem[7617] = 80'h01100a9e644e280a0969;
mem[7618] = 80'h00000000000000000000;
mem[7619] = 80'h00000000000000000000;
mem[7620] = 80'h00000000000000000000;
mem[7621] = 80'h10100000010000010010;
mem[7622] = 80'h00109400000208004500;
mem[7623] = 80'h0010002e2bb60000fffd;
mem[7624] = 80'h00100dc4c0550102c000;
mem[7625] = 80'h00100001ffabffabffab;
mem[7626] = 80'h00104989d4a229fa256b;
mem[7627] = 80'h001005076e751f14221e;
mem[7628] = 80'h01101ad0c2ef494c924f;
mem[7629] = 80'h00000000000000000000;
mem[7630] = 80'h10100000010000010010;
mem[7631] = 80'h00109400000208004500;
mem[7632] = 80'h0010002e2bb70000fffd;
mem[7633] = 80'h00100dc3c0550102c000;
mem[7634] = 80'h00100001ffabffabffab;
mem[7635] = 80'h001048f80a8ef183e7d4;
mem[7636] = 80'h0010ced5e998eac3aa4f;
mem[7637] = 80'h01107cbb08e3756ebc37;
mem[7638] = 80'h00000000000000000000;
mem[7639] = 80'h00000000000000000000;
mem[7640] = 80'h00000000000000000000;
mem[7641] = 80'h10100000010000010010;
mem[7642] = 80'h00109400000208004500;
mem[7643] = 80'h0010002e2bb80000fffd;
mem[7644] = 80'h00100dc2c0550102c000;
mem[7645] = 80'h00100001ffabffabffab;
mem[7646] = 80'h001047c05d778bd33a6a;
mem[7647] = 80'h001074d94cad66d16ad5;
mem[7648] = 80'h0110b28b4ed1c578705c;
mem[7649] = 80'h00000000000000000000;
mem[7650] = 80'h00000000000000000000;
mem[7651] = 80'h00000000000000000000;
mem[7652] = 80'h00000000000000000000;
mem[7653] = 80'h10100000010000010010;
mem[7654] = 80'h00109400000208004500;
mem[7655] = 80'h0010002e2bb90000fffd;
mem[7656] = 80'h00100dc1c0550102c000;
mem[7657] = 80'h00100001ffabffabffab;
mem[7658] = 80'h001046b1835b53aaf8d5;
mem[7659] = 80'h0010bf0bcb4093012a84;
mem[7660] = 80'h0110ce8dd31236505215;
mem[7661] = 80'h00000000000000000000;
mem[7662] = 80'h00000000000000000000;
mem[7663] = 80'h00000000000000000000;
mem[7664] = 80'h10100000010000010010;
mem[7665] = 80'h00109400000208004500;
mem[7666] = 80'h0010002e2bba0000fffd;
mem[7667] = 80'h00100dc0c0550102c000;
mem[7668] = 80'h00100001ffabffabffab;
mem[7669] = 80'h00104523e12e3b20bf15;
mem[7670] = 80'h0010e37c43768d71e876;
mem[7671] = 80'h01103cc405d84d616c11;
mem[7672] = 80'h00000000000000000000;
mem[7673] = 80'h00000000000000000000;
mem[7674] = 80'h00000000000000000000;
mem[7675] = 80'h10100000010000010010;
mem[7676] = 80'h00109400000208004500;
mem[7677] = 80'h0010002e2bbb0000fffd;
mem[7678] = 80'h00100dbfc0550102c000;
mem[7679] = 80'h00100001ffabffabffab;
mem[7680] = 80'h001044523f02e3597daa;
mem[7681] = 80'h001028aec49b78a1ab27;
mem[7682] = 80'h01101591f50254c0828e;
mem[7683] = 80'h00000000000000000000;
mem[7684] = 80'h10100000010000010010;
mem[7685] = 80'h00109400000208004500;
mem[7686] = 80'h0010002e2bbc0000fffd;
mem[7687] = 80'h00100dbec0550102c000;
mem[7688] = 80'h00100001ffabffabffab;
mem[7689] = 80'h00104376fbe8324df22a;
mem[7690] = 80'h00109041d5f7444008c2;
mem[7691] = 80'h011018e3d009c48c3699;
mem[7692] = 80'h00000000000000000000;
mem[7693] = 80'h00000000000000000000;
mem[7694] = 80'h00000000000000000000;
mem[7695] = 80'h10100000010000010010;
mem[7696] = 80'h00109400000208004500;
mem[7697] = 80'h0010002e2bbd0000fffd;
mem[7698] = 80'h00100dbdc0550102c000;
mem[7699] = 80'h00100001ffabffabffab;
mem[7700] = 80'h0010420725c4ea343095;
mem[7701] = 80'h00105b93521ab1904793;
mem[7702] = 80'h011074db61bdd606fea8;
mem[7703] = 80'h00000000000000000000;
mem[7704] = 80'h10100000010000010010;
mem[7705] = 80'h00109400000208004500;
mem[7706] = 80'h0010002e2bbe0000fffd;
mem[7707] = 80'h00100dbcc0550102c000;
mem[7708] = 80'h00100001ffabffabffab;
mem[7709] = 80'h0010419547b182be7755;
mem[7710] = 80'h001007e4da2cafe08c61;
mem[7711] = 80'h01103c0a2248b17250b0;
mem[7712] = 80'h00000000000000000000;
mem[7713] = 80'h00000000000000000000;
mem[7714] = 80'h00000000000000000000;
mem[7715] = 80'h00000000000000000000;
mem[7716] = 80'h10100000010000010010;
mem[7717] = 80'h00109400000208004500;
mem[7718] = 80'h0010002e2bbf0000fffd;
mem[7719] = 80'h00100dbbc0550102c000;
mem[7720] = 80'h00100001ffabffabffab;
mem[7721] = 80'h001040e4999d5ac7b5ea;
mem[7722] = 80'h0010cc365dc15a30f730;
mem[7723] = 80'h01109963000fce710a8e;
mem[7724] = 80'h00000000000000000000;
mem[7725] = 80'h00000000000000000000;
mem[7726] = 80'h00000000000000000000;
mem[7727] = 80'h10100000010000010010;
mem[7728] = 80'h00109400000208004500;
mem[7729] = 80'h0010002e2bc00000fffd;
mem[7730] = 80'h00100dbac0550102c000;
mem[7731] = 80'h00100001ffabffabffab;
mem[7732] = 80'h00103f733c90812c1520;
mem[7733] = 80'h00106f6ee3ecf3973257;
mem[7734] = 80'h0110ec16884e7a028c49;
mem[7735] = 80'h00000000000000000000;
mem[7736] = 80'h00000000000000000000;
mem[7737] = 80'h00000000000000000000;
mem[7738] = 80'h10100000010000010010;
mem[7739] = 80'h00109400000208004500;
mem[7740] = 80'h0010002e2bc10000fffd;
mem[7741] = 80'h00100db9c0550102c000;
mem[7742] = 80'h00100001ffabffabffab;
mem[7743] = 80'h00103e02e2bc5955d79f;
mem[7744] = 80'h0010a4bc64010646b206;
mem[7745] = 80'h0110b1743bcc04ecbdea;
mem[7746] = 80'h00000000000000000000;
mem[7747] = 80'h10100000010000010010;
mem[7748] = 80'h00109400000208004500;
mem[7749] = 80'h0010002e2bc20000fffd;
mem[7750] = 80'h00100db8c0550102c000;
mem[7751] = 80'h00100001ffabffabffab;
mem[7752] = 80'h00103d9080c931df905f;
mem[7753] = 80'h0010f8cbec37183622f4;
mem[7754] = 80'h01102be03359f8a96930;
mem[7755] = 80'h00000000000000000000;
mem[7756] = 80'h00000000000000000000;
mem[7757] = 80'h00000000000000000000;
mem[7758] = 80'h10100000010000010010;
mem[7759] = 80'h00109400000208004500;
mem[7760] = 80'h0010002e2bc30000fffd;
mem[7761] = 80'h00100db7c0550102c000;
mem[7762] = 80'h00100001ffabffabffab;
mem[7763] = 80'h00103ce15ee5e9a652e0;
mem[7764] = 80'h001033196bdaede62da5;
mem[7765] = 80'h01104a14231ed64251b5;
mem[7766] = 80'h00000000000000000000;
mem[7767] = 80'h00000000000000000000;
mem[7768] = 80'h00000000000000000000;
mem[7769] = 80'h10100000010000010010;
mem[7770] = 80'h00109400000208004500;
mem[7771] = 80'h0010002e2bc40000fffd;
mem[7772] = 80'h00100db6c0550102c000;
mem[7773] = 80'h00100001ffabffabffab;
mem[7774] = 80'h00103bc59a0f38b2dd60;
mem[7775] = 80'h00108bf67ab6d1075640;
mem[7776] = 80'h0110dbe80a3ac78ad147;
mem[7777] = 80'h00000000000000000000;
mem[7778] = 80'h10100000010000010010;
mem[7779] = 80'h00109400000208004500;
mem[7780] = 80'h0010002e2bc50000fffd;
mem[7781] = 80'h00100db5c0550102c000;
mem[7782] = 80'h00100001ffabffabffab;
mem[7783] = 80'h00103ab44423e0cb1fdf;
mem[7784] = 80'h00104024fd5b24d72f11;
mem[7785] = 80'h011018e3d631080d921c;
mem[7786] = 80'h00000000000000000000;
mem[7787] = 80'h00000000000000000000;
mem[7788] = 80'h00000000000000000000;
mem[7789] = 80'h00000000000000000000;
mem[7790] = 80'h10100000010000010010;
mem[7791] = 80'h00109400000208004500;
mem[7792] = 80'h0010002e2bc60000fffd;
mem[7793] = 80'h00100db4c0550102c000;
mem[7794] = 80'h00100001ffabffabffab;
mem[7795] = 80'h0010392626568841581f;
mem[7796] = 80'h00101c53756d3aa766e3;
mem[7797] = 80'h01102dc85f0f0766e14b;
mem[7798] = 80'h00000000000000000000;
mem[7799] = 80'h10100000010000010010;
mem[7800] = 80'h00109400000208004500;
mem[7801] = 80'h0010002e2bc70000fffd;
mem[7802] = 80'h00100db3c0550102c000;
mem[7803] = 80'h00100001ffabffabffab;
mem[7804] = 80'h00103857f87a50389aa0;
mem[7805] = 80'h0010d781f280cf772fb2;
mem[7806] = 80'h0110eb562fd150ea4fa4;
mem[7807] = 80'h00000000000000000000;
mem[7808] = 80'h00000000000000000000;
mem[7809] = 80'h00000000000000000000;
mem[7810] = 80'h00000000000000000000;
mem[7811] = 80'h10100000010000010010;
mem[7812] = 80'h00109400000208004500;
mem[7813] = 80'h0010002e2bc80000fffd;
mem[7814] = 80'h00100db2c0550102c000;
mem[7815] = 80'h00100001ffabffabffab;
mem[7816] = 80'h0010376faf832a68471e;
mem[7817] = 80'h00106d8d57b543658f28;
mem[7818] = 80'h01102e4ce169f0cf9bdb;
mem[7819] = 80'h00000000000000000000;
mem[7820] = 80'h00000000000000000000;
mem[7821] = 80'h00000000000000000000;
mem[7822] = 80'h10100000010000010010;
mem[7823] = 80'h00109400000208004500;
mem[7824] = 80'h0010002e2bc90000fffd;
mem[7825] = 80'h00100db1c0550102c000;
mem[7826] = 80'h00100001ffabffabffab;
mem[7827] = 80'h0010361e71aff21185a1;
mem[7828] = 80'h0010a65fd058b6b5ce79;
mem[7829] = 80'h0110617b831b269290b1;
mem[7830] = 80'h00000000000000000000;
mem[7831] = 80'h10100000010000010010;
mem[7832] = 80'h00109400000208004500;
mem[7833] = 80'h0010002e2bca0000fffd;
mem[7834] = 80'h00100db0c0550102c000;
mem[7835] = 80'h00100001ffabffabffab;
mem[7836] = 80'h0010358c13da9a9bc261;
mem[7837] = 80'h0010fa28586ea8c68f8b;
mem[7838] = 80'h011084a94a09f9b3b865;
mem[7839] = 80'h00000000000000000000;
mem[7840] = 80'h00000000000000000000;
mem[7841] = 80'h00000000000000000000;
mem[7842] = 80'h10100000010000010010;
mem[7843] = 80'h00109400000208004500;
mem[7844] = 80'h0010002e2bcb0000fffd;
mem[7845] = 80'h00100dafc0550102c000;
mem[7846] = 80'h00100001ffabffabffab;
mem[7847] = 80'h001034fdcdf642e200de;
mem[7848] = 80'h001031fadf835d16cfda;
mem[7849] = 80'h0110f8af822cbac31aaf;
mem[7850] = 80'h00000000000000000000;
mem[7851] = 80'h00000000000000000000;
mem[7852] = 80'h00000000000000000000;
mem[7853] = 80'h10100000010000010010;
mem[7854] = 80'h00109400000208004500;
mem[7855] = 80'h0010002e2bcc0000fffd;
mem[7856] = 80'h00100daec0550102c000;
mem[7857] = 80'h00100001ffabffabffab;
mem[7858] = 80'h001033d9091c93f68f5e;
mem[7859] = 80'h00108915ceef61f78b3f;
mem[7860] = 80'h01107cf8dd809d7e5a80;
mem[7861] = 80'h00000000000000000000;
mem[7862] = 80'h10100000010000010010;
mem[7863] = 80'h00109400000208004500;
mem[7864] = 80'h0010002e2bcd0000fffd;
mem[7865] = 80'h00100dadc0550102c000;
mem[7866] = 80'h00100001ffabffabffab;
mem[7867] = 80'h001032a8d7304b8f4de1;
mem[7868] = 80'h001042c749029427836e;
mem[7869] = 80'h0110849b34bb143061fe;
mem[7870] = 80'h00000000000000000000;
mem[7871] = 80'h00000000000000000000;
mem[7872] = 80'h00000000000000000000;
mem[7873] = 80'h00000000000000000000;
mem[7874] = 80'h10100000010000010010;
mem[7875] = 80'h00109400000208004500;
mem[7876] = 80'h0010002e2bce0000fffd;
mem[7877] = 80'h00100dacc0550102c000;
mem[7878] = 80'h00100001ffabffabffab;
mem[7879] = 80'h0010313ab54523050a21;
mem[7880] = 80'h00101eb0c1348a570a9c;
mem[7881] = 80'h0110a7e4cf9c34785fdf;
mem[7882] = 80'h00000000000000000000;
mem[7883] = 80'h00000000000000000000;
mem[7884] = 80'h00000000000000000000;
mem[7885] = 80'h10100000010000010010;
mem[7886] = 80'h00109400000208004500;
mem[7887] = 80'h0010002e2bcf0000fffd;
mem[7888] = 80'h00100dabc0550102c000;
mem[7889] = 80'h00100001ffabffabffab;
mem[7890] = 80'h0010304b6b69fb7cc89e;
mem[7891] = 80'h0010d56246d97f8793cd;
mem[7892] = 80'h0110745dfc406e62504d;
mem[7893] = 80'h00000000000000000000;
mem[7894] = 80'h10100000010000010010;
mem[7895] = 80'h00109400000208004500;
mem[7896] = 80'h0010002e2bd00000fffd;
mem[7897] = 80'h00100daac0550102c000;
mem[7898] = 80'h00100001ffabffabffab;
mem[7899] = 80'h00102f4a1ab7d7a4b15c;
mem[7900] = 80'h00106aa98b5f927269a8;
mem[7901] = 80'h01105d75dd63d946ac48;
mem[7902] = 80'h00000000000000000000;
mem[7903] = 80'h00000000000000000000;
mem[7904] = 80'h00000000000000000000;
mem[7905] = 80'h10100000010000010010;
mem[7906] = 80'h00109400000208004500;
mem[7907] = 80'h0010002e2bd10000fffd;
mem[7908] = 80'h00100da9c0550102c000;
mem[7909] = 80'h00100001ffabffabffab;
mem[7910] = 80'h00102e3bc49b0fdd73e3;
mem[7911] = 80'h0010a17b0cb267a268f9;
mem[7912] = 80'h01101f8eeb105c0ef0ee;
mem[7913] = 80'h00000000000000000000;
mem[7914] = 80'h00000000000000000000;
mem[7915] = 80'h00000000000000000000;
mem[7916] = 80'h10100000010000010010;
mem[7917] = 80'h00109400000208004500;
mem[7918] = 80'h0010002e2bd20000fffd;
mem[7919] = 80'h00100da8c0550102c000;
mem[7920] = 80'h00100001ffabffabffab;
mem[7921] = 80'h00102da9a6ee67573423;
mem[7922] = 80'h0010fd0c848479d2db0b;
mem[7923] = 80'h0110d6afe2cd6c582dce;
mem[7924] = 80'h00000000000000000000;
mem[7925] = 80'h00000000000000000000;
mem[7926] = 80'h00000000000000000000;
mem[7927] = 80'h10100000010000010010;
mem[7928] = 80'h00109400000208004500;
mem[7929] = 80'h0010002e2bd30000fffd;
mem[7930] = 80'h00100da7c0550102c000;
mem[7931] = 80'h00100001ffabffabffab;
mem[7932] = 80'h00102cd878c2bf2ef69c;
mem[7933] = 80'h001036de03698c02985a;
mem[7934] = 80'h0110fffa45fa9377144e;
mem[7935] = 80'h00000000000000000000;
mem[7936] = 80'h10100000010000010010;
mem[7937] = 80'h00109400000208004500;
mem[7938] = 80'h0010002e2bd40000fffd;
mem[7939] = 80'h00100da6c0550102c000;
mem[7940] = 80'h00100001ffabffabffab;
mem[7941] = 80'h00102bfcbc286e3a791c;
mem[7942] = 80'h00108e311205b0e22bbf;
mem[7943] = 80'h0110c6cbecdfcbb474ba;
mem[7944] = 80'h00000000000000000000;
mem[7945] = 80'h00000000000000000000;
mem[7946] = 80'h00000000000000000000;
mem[7947] = 80'h00000000000000000000;
mem[7948] = 80'h10100000010000010010;
mem[7949] = 80'h00109400000208004500;
mem[7950] = 80'h0010002e2bd50000fffd;
mem[7951] = 80'h00100da5c0550102c000;
mem[7952] = 80'h00100001ffabffabffab;
mem[7953] = 80'h00102a8d6204b643bba3;
mem[7954] = 80'h001045e395e8453274ee;
mem[7955] = 80'h0110a980c21960c3ba84;
mem[7956] = 80'h00000000000000000000;
mem[7957] = 80'h10100000010000010010;
mem[7958] = 80'h00109400000208004500;
mem[7959] = 80'h0010002e2bd60000fffd;
mem[7960] = 80'h00100da4c0550102c000;
mem[7961] = 80'h00100001ffabffabffab;
mem[7962] = 80'h0010291f0071dec9fc63;
mem[7963] = 80'h001019941dde5b42bc1c;
mem[7964] = 80'h0110b402f86dd9dbebec;
mem[7965] = 80'h00000000000000000000;
mem[7966] = 80'h00000000000000000000;
mem[7967] = 80'h00000000000000000000;
mem[7968] = 80'h00000000000000000000;
mem[7969] = 80'h10100000010000010010;
mem[7970] = 80'h00109400000208004500;
mem[7971] = 80'h0010002e2bd70000fffd;
mem[7972] = 80'h00100da3c0550102c000;
mem[7973] = 80'h00100001ffabffabffab;
mem[7974] = 80'h0010286ede5d06b03edc;
mem[7975] = 80'h0010d2469a33ae92f44d;
mem[7976] = 80'h011041ad629f462b6799;
mem[7977] = 80'h00000000000000000000;
mem[7978] = 80'h00000000000000000000;
mem[7979] = 80'h00000000000000000000;
mem[7980] = 80'h10100000010000010010;
mem[7981] = 80'h00109400000208004500;
mem[7982] = 80'h0010002e2bd80000fffd;
mem[7983] = 80'h00100da2c0550102c000;
mem[7984] = 80'h00100001ffabffabffab;
mem[7985] = 80'h0010275689a47ce0e362;
mem[7986] = 80'h0010684a3f06228035d7;
mem[7987] = 80'h0110bcac326ddc413c79;
mem[7988] = 80'h00000000000000000000;
mem[7989] = 80'h10100000010000010010;
mem[7990] = 80'h00109400000208004500;
mem[7991] = 80'h0010002e2bd90000fffd;
mem[7992] = 80'h00100da1c0550102c000;
mem[7993] = 80'h00100001ffabffabffab;
mem[7994] = 80'h001026275788a49921dd;
mem[7995] = 80'h0010a398b8ebd750b686;
mem[7996] = 80'h011083ad4dd0362979f0;
mem[7997] = 80'h00000000000000000000;
mem[7998] = 80'h00000000000000000000;
mem[7999] = 80'h00000000000000000000;
mem[8000] = 80'h00000000000000000000;
mem[8001] = 80'h10100000010000010010;
mem[8002] = 80'h00109400000208004500;
mem[8003] = 80'h0010002e2bda0000fffd;
mem[8004] = 80'h00100da0c0550102c000;
mem[8005] = 80'h00100001ffabffabffab;
mem[8006] = 80'h001025b535fdcc13661d;
mem[8007] = 80'h0010ffef30ddc9203574;
mem[8008] = 80'h01104f19f3a0a8153b1b;
mem[8009] = 80'h00000000000000000000;
mem[8010] = 80'h10100000010000010010;
mem[8011] = 80'h00109400000208004500;
mem[8012] = 80'h0010002e2bdb0000fffd;
mem[8013] = 80'h00100d9fc0550102c000;
mem[8014] = 80'h00100001ffabffabffab;
mem[8015] = 80'h001024c4ebd1146aa4a2;
mem[8016] = 80'h0010343db7303cf02a25;
mem[8017] = 80'h01102d9eb63bc97e7041;
mem[8018] = 80'h00000000000000000000;
mem[8019] = 80'h00000000000000000000;
mem[8020] = 80'h00000000000000000000;
mem[8021] = 80'h00000000000000000000;
mem[8022] = 80'h10100000010000010010;
mem[8023] = 80'h00109400000208004500;
mem[8024] = 80'h0010002e2bdc0000fffd;
mem[8025] = 80'h00100d9ec0550102c000;
mem[8026] = 80'h00100001ffabffabffab;
mem[8027] = 80'h001023e02f3bc57e2b22;
mem[8028] = 80'h00108cd2a65c001151c0;
mem[8029] = 80'h0110bc627ae0fc5efbbd;
mem[8030] = 80'h00000000000000000000;
mem[8031] = 80'h00000000000000000000;
mem[8032] = 80'h00000000000000000000;
mem[8033] = 80'h10100000010000010010;
mem[8034] = 80'h00109400000208004500;
mem[8035] = 80'h0010002e2bdd0000fffd;
mem[8036] = 80'h00100d9dc0550102c000;
mem[8037] = 80'h00100001ffabffabffab;
mem[8038] = 80'h00102291f1171d07e99d;
mem[8039] = 80'h0010470021b1f5ded891;
mem[8040] = 80'h011003faaa95b72608a7;
mem[8041] = 80'h00000000000000000000;
mem[8042] = 80'h10100000010000010010;
mem[8043] = 80'h00109400000208004500;
mem[8044] = 80'h0010002e2bde0000fffd;
mem[8045] = 80'h00100d9cc0550102c000;
mem[8046] = 80'h00100001ffabffabffab;
mem[8047] = 80'h001021039362758dae5d;
mem[8048] = 80'h00101b77a987ebae5163;
mem[8049] = 80'h011020850519a78ce519;
mem[8050] = 80'h00000000000000000000;
mem[8051] = 80'h00000000000000000000;
mem[8052] = 80'h00000000000000000000;
mem[8053] = 80'h00000000000000000000;
mem[8054] = 80'h10100000010000010010;
mem[8055] = 80'h00109400000208004500;
mem[8056] = 80'h0010002e2bdf0000fffd;
mem[8057] = 80'h00100d9bc0550102c000;
mem[8058] = 80'h00100001ffabffabffab;
mem[8059] = 80'h001020724d4eadf46ce2;
mem[8060] = 80'h0010d0a52e6a1e7e2932;
mem[8061] = 80'h0110d0bf5fe84877e6f6;
mem[8062] = 80'h00000000000000000000;
mem[8063] = 80'h10100000010000010010;
mem[8064] = 80'h00109400000208004500;
mem[8065] = 80'h0010002e2be00000fffd;
mem[8066] = 80'h00100d9ac0550102c000;
mem[8067] = 80'h00100001ffabffabffab;
mem[8068] = 80'h00101f0170de2c3d5dd8;
mem[8069] = 80'h001064e0328a304587a9;
mem[8070] = 80'h011012518460c84ab09f;
mem[8071] = 80'h00000000000000000000;
mem[8072] = 80'h00000000000000000000;
mem[8073] = 80'h00000000000000000000;
mem[8074] = 80'h00000000000000000000;
mem[8075] = 80'h10100000010000010010;
mem[8076] = 80'h00109400000208004500;
mem[8077] = 80'h0010002e2be10000fffd;
mem[8078] = 80'h00100d99c0550102c000;
mem[8079] = 80'h00100001ffabffabffab;
mem[8080] = 80'h00101e70aef2f4449f67;
mem[8081] = 80'h0010af32b567c595c7f8;
mem[8082] = 80'h01106e573e7030538d13;
mem[8083] = 80'h00000000000000000000;
mem[8084] = 80'h00000000000000000000;
mem[8085] = 80'h00000000000000000000;
mem[8086] = 80'h10100000010000010010;
mem[8087] = 80'h00109400000208004500;
mem[8088] = 80'h0010002e2be20000fffd;
mem[8089] = 80'h00100d98c0550102c000;
mem[8090] = 80'h00100001ffabffabffab;
mem[8091] = 80'h00101de2cc879cced8a7;
mem[8092] = 80'h0010f3453d51dbe5960a;
mem[8093] = 80'h0110d1a62bf17b35ab2f;
mem[8094] = 80'h00000000000000000000;
mem[8095] = 80'h10100000010000010010;
mem[8096] = 80'h00109400000208004500;
mem[8097] = 80'h0010002e2be30000fffd;
mem[8098] = 80'h00100d97c0550102c000;
mem[8099] = 80'h00100001ffabffabffab;
mem[8100] = 80'h00101c9312ab44b71a18;
mem[8101] = 80'h00103897babc2e35d75b;
mem[8102] = 80'h01109e91da7bfd3975ee;
mem[8103] = 80'h00000000000000000000;
mem[8104] = 80'h00000000000000000000;
mem[8105] = 80'h00000000000000000000;
mem[8106] = 80'h10100000010000010010;
mem[8107] = 80'h00109400000208004500;
mem[8108] = 80'h0010002e2be40000fffd;
mem[8109] = 80'h00100d96c0550102c000;
mem[8110] = 80'h00100001ffabffabffab;
mem[8111] = 80'h00101bb7d64195a39598;
mem[8112] = 80'h00108078abd012d4e2be;
mem[8113] = 80'h011021ae9f40ba43e3be;
mem[8114] = 80'h00000000000000000000;
mem[8115] = 80'h00000000000000000000;
mem[8116] = 80'h00000000000000000000;
mem[8117] = 80'h10100000010000010010;
mem[8118] = 80'h00109400000208004500;
mem[8119] = 80'h0010002e2be50000fffd;
mem[8120] = 80'h00100d95c0550102c000;
mem[8121] = 80'h00100001ffabffabffab;
mem[8122] = 80'h00101ac6086d4dda5727;
mem[8123] = 80'h00104baa2c3de7049bef;
mem[8124] = 80'h0110e2a55a49410cae90;
mem[8125] = 80'h00000000000000000000;
mem[8126] = 80'h00000000000000000000;
mem[8127] = 80'h00000000000000000000;
mem[8128] = 80'h10100000010000010010;
mem[8129] = 80'h00109400000208004500;
mem[8130] = 80'h0010002e2be60000fffd;
mem[8131] = 80'h00100d94c0550102c000;
mem[8132] = 80'h00100001ffabffabffab;
mem[8133] = 80'h001019546a18255010e7;
mem[8134] = 80'h001017dda40bf974121d;
mem[8135] = 80'h0110c1dabd0656f08e14;
mem[8136] = 80'h00000000000000000000;
mem[8137] = 80'h10100000010000010010;
mem[8138] = 80'h00109400000208004500;
mem[8139] = 80'h0010002e2be70000fffd;
mem[8140] = 80'h00100d93c0550102c000;
mem[8141] = 80'h00100001ffabffabffab;
mem[8142] = 80'h00101825b434fd29d258;
mem[8143] = 80'h0010dc0f23e60ca59b4c;
mem[8144] = 80'h01102620961b33d5cd40;
mem[8145] = 80'h00000000000000000000;
mem[8146] = 80'h00000000000000000000;
mem[8147] = 80'h00000000000000000000;
mem[8148] = 80'h10100000010000010010;
mem[8149] = 80'h00109400000208004500;
mem[8150] = 80'h0010002e2be80000fffd;
mem[8151] = 80'h00100d92c0550102c000;
mem[8152] = 80'h00100001ffabffabffab;
mem[8153] = 80'h0010171de3cd87790fe6;
mem[8154] = 80'h0010660386d380b77bd6;
mem[8155] = 80'h0110eef6955907ffa279;
mem[8156] = 80'h00000000000000000000;
mem[8157] = 80'h00000000000000000000;
mem[8158] = 80'h00000000000000000000;
mem[8159] = 80'h00000000000000000000;
mem[8160] = 80'h10100000010000010010;
mem[8161] = 80'h00109400000208004500;
mem[8162] = 80'h0010002e2be90000fffd;
mem[8163] = 80'h00100d91c0550102c000;
mem[8164] = 80'h00100001ffabffabffab;
mem[8165] = 80'h0010166c3de15f00cd59;
mem[8166] = 80'h0010add1013e75677a87;
mem[8167] = 80'h0110ac0d344c326f2f45;
mem[8168] = 80'h00000000000000000000;
mem[8169] = 80'h10100000010000010010;
mem[8170] = 80'h00109400000208004500;
mem[8171] = 80'h0010002e2bea0000fffd;
mem[8172] = 80'h00100d90c0550102c000;
mem[8173] = 80'h00100001ffabffabffab;
mem[8174] = 80'h001015fe5f94378a8a99;
mem[8175] = 80'h0010f1a689086b17fa75;
mem[8176] = 80'h011035eab222e3cf4057;
mem[8177] = 80'h00000000000000000000;
mem[8178] = 80'h00000000000000000000;
mem[8179] = 80'h00000000000000000000;
mem[8180] = 80'h10100000010000010010;
mem[8181] = 80'h00109400000208004500;
mem[8182] = 80'h0010002e2beb0000fffd;
mem[8183] = 80'h00100d8fc0550102c000;
mem[8184] = 80'h00100001ffabffabffab;
mem[8185] = 80'h0010148f81b8eff34826;
mem[8186] = 80'h00103a740ee59ec77a24;
mem[8187] = 80'h01105fb86fa064ffcaed;
mem[8188] = 80'h00000000000000000000;
mem[8189] = 80'h00000000000000000000;
mem[8190] = 80'h00000000000000000000;
mem[8191] = 80'h00000000000000000000;
end


//*********************
//MAIN CORE
//********************* 
reg [15:0] time_cnt ;    
reg [31:0] cnt ;

initial begin
    time_cnt = 'd0 ;
    cnt      = 'd0 ;
end

always @(posedge clk) begin

    if ( time_cnt == 'd1000 ) begin
        time_cnt <= time_cnt ;
    end
    else begin
        time_cnt <= time_cnt+1'b1 ;
    end
end

always @(posedge clk) begin

    if ( time_cnt >'d900 ) begin
        if ( cnt == 'd8191 ) begin
            cnt <= 'd0 ;
        end
        else begin
           cnt <= cnt+1'b1 ; 
        end
    end
    else begin
        cnt <= 'd0 ;
    end
end

wire [12:0] rd_addr ;

assign rd_addr = cnt[12:0] ;

always @(posedge clk) begin
	dout_ff <= mem[rd_addr] ;
end


assign sop  = dout_ff[76] ;
assign eop  = dout_ff[72] ;
assign dval = dout_ff[68] ;
assign mod  = dout_ff[66:64] ;
assign dout = dout_ff[63:0] ;


//*********************
endmodule   