
// **************************************************************
// COPYRIGHT(c)2015, Xidian University
// All rights reserved.
//
// IP LIB INDEX :  
// IP Name      :      
// File name    : 
// Module name  : 
// Full name    :  
//
// Author       : Liu-Huan 
// Email        : assasin9997@163.com 
// Data         : 
// Version      : V 1.0 
// 
// Abstract     : 
// Called by    :  
// 
// Modification history
// -----------------------------------------------------------------
// 
// 
//
// *****************************************************************

// *******************
// TIMESCALE
// ******************* 
`timescale 1ns/1ps 

// *******************
// INFORMATION
// *******************


//*******************
//DEFINE(s)
//*******************
//`define UDLY 1    //Unit delay, for non-blocking assignments in sequential logic


//*******************
//DEFINE MODULE PORT
//*******************
module  data_source_random   (     
            input 				clk     ,
            output  			sop     ,
            output  			eop     ,
            output  			dval    ,
            output  [2:0] 		mod     ,
            output  [63:0] 		dout         
              ) ;

//*******************
//DEFINE LOCAL PARAMETER
//*******************
//parameter(s)
                                    
 

//*********************
//INNER SIGNAL DECLARATION
//*********************
//REGS
  reg [79:0] mem [0:8191] ;
  reg [79:0] dout_ff = 80'b0 ;

//WIRES
 

//*********************
//INSTANTCE MODULE
//*********************

initial begin
mem[0]    = 80'h00000000000000000000;
mem[1]    = 80'h10100000010000010010;
mem[2]    = 80'h00109400000208004500;
mem[3]    = 80'h0010028f899a0000fffd;
mem[4]    = 80'h0010ad7ec0550102c000;
mem[5]    = 80'h00100001ffabffabffab;
mem[6]    = 80'h0010ffabffabffabffab;
mem[7]    = 80'h0010ffabffabffabffab;
mem[8]    = 80'h0010ffabffabffabffab;
mem[9]    = 80'h0010ffabffabffabffab;
mem[10]   = 80'h0010ffabffabffabffab;
mem[11]   = 80'h0010ffabffabffabffab;
mem[12]   = 80'h0010ffabffabffabffab;
mem[13]   = 80'h0010ffabffabffabffab;
mem[14]   = 80'h0010ffabffabffabffab;
mem[15]   = 80'h0010ffabffabffabffab;
mem[16]   = 80'h0010ffabffabffabffab;
mem[17]   = 80'h0010ffabffabffabffab;
mem[18]   = 80'h0010ffabffabffabffab;
mem[19]   = 80'h0010ffabffabffabffab;
mem[20]   = 80'h0010ffabffabffabffab;
mem[21]   = 80'h0010ffabffabffabffab;
mem[22]   = 80'h0010ffabffabffabffab;
mem[23]   = 80'h0010ffabffabffabffab;
mem[24]   = 80'h0010ffabffabffabffab;
mem[25]   = 80'h0010ffabffabffabffab;
mem[26]   = 80'h0010ffabffabffabffab;
mem[27]   = 80'h0010ffabffabffabffab;
mem[28]   = 80'h0010ffabffabffabffab;
mem[29]   = 80'h0010ffabffabffabffab;
mem[30]   = 80'h0010ffabffabffabffab;
mem[31]   = 80'h0010ffabffabffabffab;
mem[32]   = 80'h0010ffabffabffabffab;
mem[33]   = 80'h0010ffabffabffabffab;
mem[34]   = 80'h0010ffabffabffabffab;
mem[35]   = 80'h0010ffabffabffabffab;
mem[36]   = 80'h0010ffabffabffabffab;
mem[37]   = 80'h0010ffabffabffabffab;
mem[38]   = 80'h0010ffabffabffabffab;
mem[39]   = 80'h0010ffabffabffabffab;
mem[40]   = 80'h0010ffabffabffabffab;
mem[41]   = 80'h0010ffabffabffabffab;
mem[42]   = 80'h0010ffabffabffabffab;
mem[43]   = 80'h0010ffabffabffabffab;
mem[44]   = 80'h0010ffabffabffabffab;
mem[45]   = 80'h0010ffabffabffabffab;
mem[46]   = 80'h0010ffabffabffabffab;
mem[47]   = 80'h0010ffabffabffabffab;
mem[48]   = 80'h0010ffabffabffabffab;
mem[49]   = 80'h0010ffabffabffabffab;
mem[50]   = 80'h0010ffabffabffabffab;
mem[51]   = 80'h0010ffabffabffabffab;
mem[52]   = 80'h0010ffabffabffabffab;
mem[53]   = 80'h0010ffabffabffabffab;
mem[54]   = 80'h0010ffabffabffabffab;
mem[55]   = 80'h0010ffabffabffabffab;
mem[56]   = 80'h0010ffabffabffabffab;
mem[57]   = 80'h0010ffabffabffabffab;
mem[58]   = 80'h0010ffabffabffabffab;
mem[59]   = 80'h0010ffabffabffabffab;
mem[60]   = 80'h0010ffabffabffabffab;
mem[61]   = 80'h0010ffabffabffabffab;
mem[62]   = 80'h0010ffabffabffabffab;
mem[63]   = 80'h0010ffabffabffabffab;
mem[64]   = 80'h0010ffabffabffabffab;
mem[65]   = 80'h0010ffabffabffabffab;
mem[66]   = 80'h0010ffabffabffabffab;
mem[67]   = 80'h0010ffabffabffabffab;
mem[68]   = 80'h0010ffabffabffabffab;
mem[69]   = 80'h0010ffabffabffabffab;
mem[70]   = 80'h0010ffabffabffabffab;
mem[71]   = 80'h0010ffabffabffabffab;
mem[72]   = 80'h0010ffabffabffabffab;
mem[73]   = 80'h0010ffabffabffabffab;
mem[74]   = 80'h0010ffabffabffabffab;
mem[75]   = 80'h0010ffabffabffabffab;
mem[76]   = 80'h0010ffabffabffabffab;
mem[77]   = 80'h0010ffabffabffabffab;
mem[78]   = 80'h0010ffabffabffabffab;
mem[79]   = 80'h0010ffabffabffabffab;
mem[80]   = 80'h0010ffabffabffabffab;
mem[81]   = 80'h0010ffabffabffabffab;
mem[82]   = 80'h0010ff6551ad60965d5b;
mem[83]   = 80'h001081445092d97f0a64;
mem[84]   = 80'h00102c32d20e3c39da44;
mem[85]   = 80'h0111ec00000000000000;
mem[86]   = 80'h10100000010000010010;
mem[87]   = 80'h00109400000208004500;
mem[88]   = 80'h00100437899b0000fffd;
mem[89]   = 80'h0010abd5c0550102c000;
mem[90]   = 80'h00100001ffabffabffab;
mem[91]   = 80'h0010ffabffabffabffab;
mem[92]   = 80'h0010ffabffabffabffab;
mem[93]   = 80'h0010ffabffabffabffab;
mem[94]   = 80'h0010ffabffabffabffab;
mem[95]   = 80'h0010ffabffabffabffab;
mem[96]   = 80'h0010ffabffabffabffab;
mem[97]   = 80'h0010ffabffabffabffab;
mem[98]   = 80'h0010ffabffabffabffab;
mem[99]   = 80'h0010ffabffabffabffab;
mem[100]  = 80'h0010ffabffabffabffab;
mem[101]  = 80'h0010ffabffabffabffab;
mem[102]  = 80'h0010ffabffabffabffab;
mem[103]  = 80'h0010ffabffabffabffab;
mem[104]  = 80'h0010ffabffabffabffab;
mem[105]  = 80'h0010ffabffabffabffab;
mem[106]  = 80'h0010ffabffabffabffab;
mem[107]  = 80'h0010ffabffabffabffab;
mem[108]  = 80'h0010ffabffabffabffab;
mem[109]  = 80'h0010ffabffabffabffab;
mem[110]  = 80'h0010ffabffabffabffab;
mem[111]  = 80'h0010ffabffabffabffab;
mem[112]  = 80'h0010ffabffabffabffab;
mem[113]  = 80'h0010ffabffabffabffab;
mem[114]  = 80'h0010ffabffabffabffab;
mem[115]  = 80'h0010ffabffabffabffab;
mem[116]  = 80'h0010ffabffabffabffab;
mem[117]  = 80'h0010ffabffabffabffab;
mem[118]  = 80'h0010ffabffabffabffab;
mem[119]  = 80'h0010ffabffabffabffab;
mem[120]  = 80'h0010ffabffabffabffab;
mem[121]  = 80'h0010ffabffabffabffab;
mem[122]  = 80'h0010ffabffabffabffab;
mem[123]  = 80'h0010ffabffabffabffab;
mem[124]  = 80'h0010ffabffabffabffab;
mem[125]  = 80'h0010ffabffabffabffab;
mem[126]  = 80'h0010ffabffabffabffab;
mem[127]  = 80'h0010ffabffabffabffab;
mem[128]  = 80'h0010ffabffabffabffab;
mem[129]  = 80'h0010ffabffabffabffab;
mem[130]  = 80'h0010ffabffabffabffab;
mem[131]  = 80'h0010ffabffabffabffab;
mem[132]  = 80'h0010ffabffabffabffab;
mem[133]  = 80'h0010ffabffabffabffab;
mem[134]  = 80'h0010ffabffabffabffab;
mem[135]  = 80'h0010ffabffabffabffab;
mem[136]  = 80'h0010ffabffabffabffab;
mem[137]  = 80'h0010ffabffabffabffab;
mem[138]  = 80'h0010ffabffabffabffab;
mem[139]  = 80'h0010ffabffabffabffab;
mem[140]  = 80'h0010ffabffabffabffab;
mem[141]  = 80'h0010ffabffabffabffab;
mem[142]  = 80'h0010ffabffabffabffab;
mem[143]  = 80'h0010ffabffabffabffab;
mem[144]  = 80'h0010ffabffabffabffab;
mem[145]  = 80'h0010ffabffabffabffab;
mem[146]  = 80'h0010ffabffabffabffab;
mem[147]  = 80'h0010ffabffabffabffab;
mem[148]  = 80'h0010ffabffabffabffab;
mem[149]  = 80'h0010ffabffabffabffab;
mem[150]  = 80'h0010ffabffabffabffab;
mem[151]  = 80'h0010ffabffabffabffab;
mem[152]  = 80'h0010ffabffabffabffab;
mem[153]  = 80'h0010ffabffabffabffab;
mem[154]  = 80'h0010ffabffabffabffab;
mem[155]  = 80'h0010ffabffabffabffab;
mem[156]  = 80'h0010ffabffabffabffab;
mem[157]  = 80'h0010ffabffabffabffab;
mem[158]  = 80'h0010ffabffabffabffab;
mem[159]  = 80'h0010ffabffabffabffab;
mem[160]  = 80'h0010ffabffabffabffab;
mem[161]  = 80'h0010ffabffabffabffab;
mem[162]  = 80'h0010ffabffabffabffab;
mem[163]  = 80'h0010ffabffabffabffab;
mem[164]  = 80'h0010ffabffabffabffab;
mem[165]  = 80'h0010ffabffabffabffab;
mem[166]  = 80'h0010ffabffabffabffab;
mem[167]  = 80'h0010ffabffabffabffab;
mem[168]  = 80'h0010ffabffabffabffab;
mem[169]  = 80'h0010ffabffabffabffab;
mem[170]  = 80'h0010ffabffabffabffab;
mem[171]  = 80'h0010ffabffabffabffab;
mem[172]  = 80'h0010ffabffabffabffab;
mem[173]  = 80'h0010ffabffabffabffab;
mem[174]  = 80'h0010ffabffabffabffab;
mem[175]  = 80'h0010ffabffabffabffab;
mem[176]  = 80'h0010ffabffabffabffab;
mem[177]  = 80'h0010ffabffabffabffab;
mem[178]  = 80'h0010ffabffabffabffab;
mem[179]  = 80'h0010ffabffabffabffab;
mem[180]  = 80'h0010ffabffabffabffab;
mem[181]  = 80'h0010ffabffabffabffab;
mem[182]  = 80'h0010ffabffabffabffab;
mem[183]  = 80'h0010ffabffabffabffab;
mem[184]  = 80'h0010ffabffabffabffab;
mem[185]  = 80'h0010ffabffabffabffab;
mem[186]  = 80'h0010ffabffabffabffab;
mem[187]  = 80'h0010ffabffabffabffab;
mem[188]  = 80'h0010ffabffabffabffab;
mem[189]  = 80'h0010ffabffabffabffab;
mem[190]  = 80'h0010ffabffabffabffab;
mem[191]  = 80'h0010ffabffabffabffab;
mem[192]  = 80'h0010ffabffabffabffab;
mem[193]  = 80'h0010ffabffabffabffab;
mem[194]  = 80'h0010ffabffabffabffab;
mem[195]  = 80'h0010ffabffabffabffab;
mem[196]  = 80'h0010ffabffabffabffab;
mem[197]  = 80'h0010ffabffabffabffab;
mem[198]  = 80'h0010ffabffabffabffab;
mem[199]  = 80'h0010ffabffabffabffab;
mem[200]  = 80'h0010ffabffabffabffab;
mem[201]  = 80'h0010ffabffabffabffab;
mem[202]  = 80'h0010ffabffabffabffab;
mem[203]  = 80'h0010ffabffabffabffab;
mem[204]  = 80'h0010ffabffabffabffab;
mem[205]  = 80'h0010ffabffabffabffab;
mem[206]  = 80'h0010ffabffabffabffab;
mem[207]  = 80'h0010ffabffabffabffab;
mem[208]  = 80'h0010ffabffabffabffab;
mem[209]  = 80'h0010ffabffabffabffab;
mem[210]  = 80'h0010ffabffabffabffab;
mem[211]  = 80'h0010ffabffabffabffab;
mem[212]  = 80'h0010ffabffabffabffab;
mem[213]  = 80'h0010ffabffabffabffab;
mem[214]  = 80'h0010ffabffabffabffab;
mem[215]  = 80'h0010ffabffabffabffab;
mem[216]  = 80'h0010ffabffabffabffab;
mem[217]  = 80'h0010ffabffabffabffab;
mem[218]  = 80'h0010ffabffabffabffab;
mem[219]  = 80'h0010ffabffabffabffab;
mem[220]  = 80'h0010ff6420734c4e2499;
mem[221]  = 80'h00103e8f8215348ad960;
mem[222]  = 80'h00107dd68cda9563f9a7;
mem[223]  = 80'h01118200000000000000;
mem[224]  = 80'h00000000000000000000;
mem[225]  = 80'h00000000000000000000;
mem[226]  = 80'h00000000000000000000;
mem[227]  = 80'h00000000000000000000;
mem[228]  = 80'h00000000000000000000;
mem[229]  = 80'h00000000000000000000;
mem[230]  = 80'h00000000000000000000;
mem[231]  = 80'h00000000000000000000;
mem[232]  = 80'h00000000000000000000;
mem[233]  = 80'h10100000010000010010;
mem[234]  = 80'h00109400000208004500;
mem[235]  = 80'h0010050a899c0000fffd;
mem[236]  = 80'h0010ab01c0550102c000;
mem[237]  = 80'h00100001ffabffabffab;
mem[238]  = 80'h0010ffabffabffabffab;
mem[239]  = 80'h0010ffabffabffabffab;
mem[240]  = 80'h0010ffabffabffabffab;
mem[241]  = 80'h0010ffabffabffabffab;
mem[242]  = 80'h0010ffabffabffabffab;
mem[243]  = 80'h0010ffabffabffabffab;
mem[244]  = 80'h0010ffabffabffabffab;
mem[245]  = 80'h0010ffabffabffabffab;
mem[246]  = 80'h0010ffabffabffabffab;
mem[247]  = 80'h0010ffabffabffabffab;
mem[248]  = 80'h0010ffabffabffabffab;
mem[249]  = 80'h0010ffabffabffabffab;
mem[250]  = 80'h0010ffabffabffabffab;
mem[251]  = 80'h0010ffabffabffabffab;
mem[252]  = 80'h0010ffabffabffabffab;
mem[253]  = 80'h0010ffabffabffabffab;
mem[254]  = 80'h0010ffabffabffabffab;
mem[255]  = 80'h0010ffabffabffabffab;
mem[256]  = 80'h0010ffabffabffabffab;
mem[257]  = 80'h0010ffabffabffabffab;
mem[258]  = 80'h0010ffabffabffabffab;
mem[259]  = 80'h0010ffabffabffabffab;
mem[260]  = 80'h0010ffabffabffabffab;
mem[261]  = 80'h0010ffabffabffabffab;
mem[262]  = 80'h0010ffabffabffabffab;
mem[263]  = 80'h0010ffabffabffabffab;
mem[264]  = 80'h0010ffabffabffabffab;
mem[265]  = 80'h0010ffabffabffabffab;
mem[266]  = 80'h0010ffabffabffabffab;
mem[267]  = 80'h0010ffabffabffabffab;
mem[268]  = 80'h0010ffabffabffabffab;
mem[269]  = 80'h0010ffabffabffabffab;
mem[270]  = 80'h0010ffabffabffabffab;
mem[271]  = 80'h0010ffabffabffabffab;
mem[272]  = 80'h0010ffabffabffabffab;
mem[273]  = 80'h0010ffabffabffabffab;
mem[274]  = 80'h0010ffabffabffabffab;
mem[275]  = 80'h0010ffabffabffabffab;
mem[276]  = 80'h0010ffabffabffabffab;
mem[277]  = 80'h0010ffabffabffabffab;
mem[278]  = 80'h0010ffabffabffabffab;
mem[279]  = 80'h0010ffabffabffabffab;
mem[280]  = 80'h0010ffabffabffabffab;
mem[281]  = 80'h0010ffabffabffabffab;
mem[282]  = 80'h0010ffabffabffabffab;
mem[283]  = 80'h0010ffabffabffabffab;
mem[284]  = 80'h0010ffabffabffabffab;
mem[285]  = 80'h0010ffabffabffabffab;
mem[286]  = 80'h0010ffabffabffabffab;
mem[287]  = 80'h0010ffabffabffabffab;
mem[288]  = 80'h0010ffabffabffabffab;
mem[289]  = 80'h0010ffabffabffabffab;
mem[290]  = 80'h0010ffabffabffabffab;
mem[291]  = 80'h0010ffabffabffabffab;
mem[292]  = 80'h0010ffabffabffabffab;
mem[293]  = 80'h0010ffabffabffabffab;
mem[294]  = 80'h0010ffabffabffabffab;
mem[295]  = 80'h0010ffabffabffabffab;
mem[296]  = 80'h0010ffabffabffabffab;
mem[297]  = 80'h0010ffabffabffabffab;
mem[298]  = 80'h0010ffabffabffabffab;
mem[299]  = 80'h0010ffabffabffabffab;
mem[300]  = 80'h0010ffabffabffabffab;
mem[301]  = 80'h0010ffabffabffabffab;
mem[302]  = 80'h0010ffabffabffabffab;
mem[303]  = 80'h0010ffabffabffabffab;
mem[304]  = 80'h0010ffabffabffabffab;
mem[305]  = 80'h0010ffabffabffabffab;
mem[306]  = 80'h0010ffabffabffabffab;
mem[307]  = 80'h0010ffabffabffabffab;
mem[308]  = 80'h0010ffabffabffabffab;
mem[309]  = 80'h0010ffabffabffabffab;
mem[310]  = 80'h0010ffabffabffabffab;
mem[311]  = 80'h0010ffabffabffabffab;
mem[312]  = 80'h0010ffabffabffabffab;
mem[313]  = 80'h0010ffabffabffabffab;
mem[314]  = 80'h0010ffabffabffabffab;
mem[315]  = 80'h0010ffabffabffabffab;
mem[316]  = 80'h0010ffabffabffabffab;
mem[317]  = 80'h0010ffabffabffabffab;
mem[318]  = 80'h0010ffabffabffabffab;
mem[319]  = 80'h0010ffabffabffabffab;
mem[320]  = 80'h0010ffabffabffabffab;
mem[321]  = 80'h0010ffabffabffabffab;
mem[322]  = 80'h0010ffabffabffabffab;
mem[323]  = 80'h0010ffabffabffabffab;
mem[324]  = 80'h0010ffabffabffabffab;
mem[325]  = 80'h0010ffabffabffabffab;
mem[326]  = 80'h0010ffabffabffabffab;
mem[327]  = 80'h0010ffabffabffabffab;
mem[328]  = 80'h0010ffabffabffabffab;
mem[329]  = 80'h0010ffabffabffabffab;
mem[330]  = 80'h0010ffabffabffabffab;
mem[331]  = 80'h0010ffabffabffabffab;
mem[332]  = 80'h0010ffabffabffabffab;
mem[333]  = 80'h0010ffabffabffabffab;
mem[334]  = 80'h0010ffabffabffabffab;
mem[335]  = 80'h0010ffabffabffabffab;
mem[336]  = 80'h0010ffabffabffabffab;
mem[337]  = 80'h0010ffabffabffabffab;
mem[338]  = 80'h0010ffabffabffabffab;
mem[339]  = 80'h0010ffabffabffabffab;
mem[340]  = 80'h0010ffabffabffabffab;
mem[341]  = 80'h0010ffabffabffabffab;
mem[342]  = 80'h0010ffabffabffabffab;
mem[343]  = 80'h0010ffabffabffabffab;
mem[344]  = 80'h0010ffabffabffabffab;
mem[345]  = 80'h0010ffabffabffabffab;
mem[346]  = 80'h0010ffabffabffabffab;
mem[347]  = 80'h0010ffabffabffabffab;
mem[348]  = 80'h0010ffabffabffabffab;
mem[349]  = 80'h0010ffabffabffabffab;
mem[350]  = 80'h0010ffabffabffabffab;
mem[351]  = 80'h0010ffabffabffabffab;
mem[352]  = 80'h0010ffabffabffabffab;
mem[353]  = 80'h0010ffabffabffabffab;
mem[354]  = 80'h0010ffabffabffabffab;
mem[355]  = 80'h0010ffabffabffabffab;
mem[356]  = 80'h0010ffabffabffabffab;
mem[357]  = 80'h0010ffabffabffabffab;
mem[358]  = 80'h0010ffabffabffabffab;
mem[359]  = 80'h0010ffabffabffabffab;
mem[360]  = 80'h0010ffabffabffabffab;
mem[361]  = 80'h0010ffabffabffabffab;
mem[362]  = 80'h0010ffabffabffabffab;
mem[363]  = 80'h0010ffabffabffabffab;
mem[364]  = 80'h0010ffabffabffabffab;
mem[365]  = 80'h0010ffabffabffabffab;
mem[366]  = 80'h0010ffabffabffabffab;
mem[367]  = 80'h0010ffabffabffabffab;
mem[368]  = 80'h0010ffabffabffabffab;
mem[369]  = 80'h0010ffabffabffabffab;
mem[370]  = 80'h0010ffabffabffabffab;
mem[371]  = 80'h0010ffabffabffabffab;
mem[372]  = 80'h0010ffabffabffabffab;
mem[373]  = 80'h0010ffabffabffabffab;
mem[374]  = 80'h0010ffabffabffabffab;
mem[375]  = 80'h0010ffabffabffabffab;
mem[376]  = 80'h0010ffabffabffabffab;
mem[377]  = 80'h0010ffabffabffabffab;
mem[378]  = 80'h0010ffabffabffabffab;
mem[379]  = 80'h0010ffabffabffabffab;
mem[380]  = 80'h0010ffabffabffabffab;
mem[381]  = 80'h0010ffabffabffabffab;
mem[382]  = 80'h0010ffabffabffabffab;
mem[383]  = 80'h0010ffabffabffabffab;
mem[384]  = 80'h0010ffabffabffabffab;
mem[385]  = 80'h0010ffabffabffabffab;
mem[386]  = 80'h0010ffabffabffabffab;
mem[387]  = 80'h0010ffabffabffabffab;
mem[388]  = 80'h0010ffabffabffabffab;
mem[389]  = 80'h0010ffabffabffabffab;
mem[390]  = 80'h0010ffabffabffabffab;
mem[391]  = 80'h0010ffabffabffabffab;
mem[392]  = 80'h0010ffabffabffabffab;
mem[393]  = 80'h0010ffabffab6304b7a6;
mem[394]  = 80'h00109f3016be376d0458;
mem[395]  = 80'h0010b63e8598ce34e994;
mem[396]  = 80'h011479b15cb800000000;
mem[397]  = 80'h00000000000000000000;
mem[398]  = 80'h00000000000000000000;
mem[399]  = 80'h00000000000000000000;
mem[400]  = 80'h00000000000000000000;
mem[401]  = 80'h00000000000000000000;
mem[402]  = 80'h00000000000000000000;
mem[403]  = 80'h00000000000000000000;
mem[404]  = 80'h00000000000000000000;
mem[405]  = 80'h00000000000000000000;
mem[406]  = 80'h00000000000000000000;
mem[407]  = 80'h00000000000000000000;
mem[408]  = 80'h00000000000000000000;
mem[409]  = 80'h00000000000000000000;
mem[410]  = 80'h00000000000000000000;
mem[411]  = 80'h00000000000000000000;
mem[412]  = 80'h10100000010000010010;
mem[413]  = 80'h00109400000208004500;
mem[414]  = 80'h00100573899d0000fffd;
mem[415]  = 80'h0010aa97c0550102c000;
mem[416]  = 80'h00100001ffabffabffab;
mem[417]  = 80'h0010ffabffabffabffab;
mem[418]  = 80'h0010ffabffabffabffab;
mem[419]  = 80'h0010ffabffabffabffab;
mem[420]  = 80'h0010ffabffabffabffab;
mem[421]  = 80'h0010ffabffabffabffab;
mem[422]  = 80'h0010ffabffabffabffab;
mem[423]  = 80'h0010ffabffabffabffab;
mem[424]  = 80'h0010ffabffabffabffab;
mem[425]  = 80'h0010ffabffabffabffab;
mem[426]  = 80'h0010ffabffabffabffab;
mem[427]  = 80'h0010ffabffabffabffab;
mem[428]  = 80'h0010ffabffabffabffab;
mem[429]  = 80'h0010ffabffabffabffab;
mem[430]  = 80'h0010ffabffabffabffab;
mem[431]  = 80'h0010ffabffabffabffab;
mem[432]  = 80'h0010ffabffabffabffab;
mem[433]  = 80'h0010ffabffabffabffab;
mem[434]  = 80'h0010ffabffabffabffab;
mem[435]  = 80'h0010ffabffabffabffab;
mem[436]  = 80'h0010ffabffabffabffab;
mem[437]  = 80'h0010ffabffabffabffab;
mem[438]  = 80'h0010ffabffabffabffab;
mem[439]  = 80'h0010ffabffabffabffab;
mem[440]  = 80'h0010ffabffabffabffab;
mem[441]  = 80'h0010ffabffabffabffab;
mem[442]  = 80'h0010ffabffabffabffab;
mem[443]  = 80'h0010ffabffabffabffab;
mem[444]  = 80'h0010ffabffabffabffab;
mem[445]  = 80'h0010ffabffabffabffab;
mem[446]  = 80'h0010ffabffabffabffab;
mem[447]  = 80'h0010ffabffabffabffab;
mem[448]  = 80'h0010ffabffabffabffab;
mem[449]  = 80'h0010ffabffabffabffab;
mem[450]  = 80'h0010ffabffabffabffab;
mem[451]  = 80'h0010ffabffabffabffab;
mem[452]  = 80'h0010ffabffabffabffab;
mem[453]  = 80'h0010ffabffabffabffab;
mem[454]  = 80'h0010ffabffabffabffab;
mem[455]  = 80'h0010ffabffabffabffab;
mem[456]  = 80'h0010ffabffabffabffab;
mem[457]  = 80'h0010ffabffabffabffab;
mem[458]  = 80'h0010ffabffabffabffab;
mem[459]  = 80'h0010ffabffabffabffab;
mem[460]  = 80'h0010ffabffabffabffab;
mem[461]  = 80'h0010ffabffabffabffab;
mem[462]  = 80'h0010ffabffabffabffab;
mem[463]  = 80'h0010ffabffabffabffab;
mem[464]  = 80'h0010ffabffabffabffab;
mem[465]  = 80'h0010ffabffabffabffab;
mem[466]  = 80'h0010ffabffabffabffab;
mem[467]  = 80'h0010ffabffabffabffab;
mem[468]  = 80'h0010ffabffabffabffab;
mem[469]  = 80'h0010ffabffabffabffab;
mem[470]  = 80'h0010ffabffabffabffab;
mem[471]  = 80'h0010ffabffabffabffab;
mem[472]  = 80'h0010ffabffabffabffab;
mem[473]  = 80'h0010ffabffabffabffab;
mem[474]  = 80'h0010ffabffabffabffab;
mem[475]  = 80'h0010ffabffabffabffab;
mem[476]  = 80'h0010ffabffabffabffab;
mem[477]  = 80'h0010ffabffabffabffab;
mem[478]  = 80'h0010ffabffabffabffab;
mem[479]  = 80'h0010ffabffabffabffab;
mem[480]  = 80'h0010ffabffabffabffab;
mem[481]  = 80'h0010ffabffabffabffab;
mem[482]  = 80'h0010ffabffabffabffab;
mem[483]  = 80'h0010ffabffabffabffab;
mem[484]  = 80'h0010ffabffabffabffab;
mem[485]  = 80'h0010ffabffabffabffab;
mem[486]  = 80'h0010ffabffabffabffab;
mem[487]  = 80'h0010ffabffabffabffab;
mem[488]  = 80'h0010ffabffabffabffab;
mem[489]  = 80'h0010ffabffabffabffab;
mem[490]  = 80'h0010ffabffabffabffab;
mem[491]  = 80'h0010ffabffabffabffab;
mem[492]  = 80'h0010ffabffabffabffab;
mem[493]  = 80'h0010ffabffabffabffab;
mem[494]  = 80'h0010ffabffabffabffab;
mem[495]  = 80'h0010ffabffabffabffab;
mem[496]  = 80'h0010ffabffabffabffab;
mem[497]  = 80'h0010ffabffabffabffab;
mem[498]  = 80'h0010ffabffabffabffab;
mem[499]  = 80'h0010ffabffabffabffab;
mem[500]  = 80'h0010ffabffabffabffab;
mem[501]  = 80'h0010ffabffabffabffab;
mem[502]  = 80'h0010ffabffabffabffab;
mem[503]  = 80'h0010ffabffabffabffab;
mem[504]  = 80'h0010ffabffabffabffab;
mem[505]  = 80'h0010ffabffabffabffab;
mem[506]  = 80'h0010ffabffabffabffab;
mem[507]  = 80'h0010ffabffabffabffab;
mem[508]  = 80'h0010ffabffabffabffab;
mem[509]  = 80'h0010ffabffabffabffab;
mem[510]  = 80'h0010ffabffabffabffab;
mem[511]  = 80'h0010ffabffabffabffab;
mem[512]  = 80'h0010ffabffabffabffab;
mem[513]  = 80'h0010ffabffabffabffab;
mem[514]  = 80'h0010ffabffabffabffab;
mem[515]  = 80'h0010ffabffabffabffab;
mem[516]  = 80'h0010ffabffabffabffab;
mem[517]  = 80'h0010ffabffabffabffab;
mem[518]  = 80'h0010ffabffabffabffab;
mem[519]  = 80'h0010ffabffabffabffab;
mem[520]  = 80'h0010ffabffabffabffab;
mem[521]  = 80'h0010ffabffabffabffab;
mem[522]  = 80'h0010ffabffabffabffab;
mem[523]  = 80'h0010ffabffabffabffab;
mem[524]  = 80'h0010ffabffabffabffab;
mem[525]  = 80'h0010ffabffabffabffab;
mem[526]  = 80'h0010ffabffabffabffab;
mem[527]  = 80'h0010ffabffabffabffab;
mem[528]  = 80'h0010ffabffabffabffab;
mem[529]  = 80'h0010ffabffabffabffab;
mem[530]  = 80'h0010ffabffabffabffab;
mem[531]  = 80'h0010ffabffabffabffab;
mem[532]  = 80'h0010ffabffabffabffab;
mem[533]  = 80'h0010ffabffabffabffab;
mem[534]  = 80'h0010ffabffabffabffab;
mem[535]  = 80'h0010ffabffabffabffab;
mem[536]  = 80'h0010ffabffabffabffab;
mem[537]  = 80'h0010ffabffabffabffab;
mem[538]  = 80'h0010ffabffabffabffab;
mem[539]  = 80'h0010ffabffabffabffab;
mem[540]  = 80'h0010ffabffabffabffab;
mem[541]  = 80'h0010ffabffabffabffab;
mem[542]  = 80'h0010ffabffabffabffab;
mem[543]  = 80'h0010ffabffabffabffab;
mem[544]  = 80'h0010ffabffabffabffab;
mem[545]  = 80'h0010ffabffabffabffab;
mem[546]  = 80'h0010ffabffabffabffab;
mem[547]  = 80'h0010ffabffabffabffab;
mem[548]  = 80'h0010ffabffabffabffab;
mem[549]  = 80'h0010ffabffabffabffab;
mem[550]  = 80'h0010ffabffabffabffab;
mem[551]  = 80'h0010ffabffabffabffab;
mem[552]  = 80'h0010ffabffabffabffab;
mem[553]  = 80'h0010ffabffabffabffab;
mem[554]  = 80'h0010ffabffabffabffab;
mem[555]  = 80'h0010ffabffabffabffab;
mem[556]  = 80'h0010ffabffabffabffab;
mem[557]  = 80'h0010ffabffabffabffab;
mem[558]  = 80'h0010ffabffabffabffab;
mem[559]  = 80'h0010ffabffabffabffab;
mem[560]  = 80'h0010ffabffabffabffab;
mem[561]  = 80'h0010ffabffabffabffab;
mem[562]  = 80'h0010ffabffabffabffab;
mem[563]  = 80'h0010ffabffabffabffab;
mem[564]  = 80'h0010ffabffabffabffab;
mem[565]  = 80'h0010ffabffabffabffab;
mem[566]  = 80'h0010ffabffabffabffab;
mem[567]  = 80'h0010ffabffabffabffab;
mem[568]  = 80'h0010ffabffabffabffab;
mem[569]  = 80'h0010ffabffabffabffab;
mem[570]  = 80'h0010ffabffabffabffab;
mem[571]  = 80'h0010ffabffabffabffab;
mem[572]  = 80'h0010ffabffabffabffab;
mem[573]  = 80'h0010ffabffabffabffab;
mem[574]  = 80'h0010ffabffabffabffab;
mem[575]  = 80'h0010ffabffabffabffab;
mem[576]  = 80'h0010ffabffabffabffab;
mem[577]  = 80'h0010ffabffabffabffab;
mem[578]  = 80'h0010ffabffabffabffab;
mem[579]  = 80'h0010ffabffabffabffab;
mem[580]  = 80'h0010ffabffabffabffab;
mem[581]  = 80'h0010ffabffabffabffab;
mem[582]  = 80'h0010ffabffabffabffab;
mem[583]  = 80'h0010ffabffabffabffab;
mem[584]  = 80'h0010ffabffabffabffab;
mem[585]  = 80'h0010ffabffabff627569;
mem[586]  = 80'h00108a4749d401fcbf83;
mem[587]  = 80'h0010b543ef4bc9bd954a;
mem[588]  = 80'h0115f1f6b98c09000000;
mem[589]  = 80'h10100000010000010010;
mem[590]  = 80'h00109400000208004500;
mem[591]  = 80'h001002d0899e0000fffd;
mem[592]  = 80'h0010ad39c0550102c000;
mem[593]  = 80'h00100001ffabffabffab;
mem[594]  = 80'h0010ffabffabffabffab;
mem[595]  = 80'h0010ffabffabffabffab;
mem[596]  = 80'h0010ffabffabffabffab;
mem[597]  = 80'h0010ffabffabffabffab;
mem[598]  = 80'h0010ffabffabffabffab;
mem[599]  = 80'h0010ffabffabffabffab;
mem[600]  = 80'h0010ffabffabffabffab;
mem[601]  = 80'h0010ffabffabffabffab;
mem[602]  = 80'h0010ffabffabffabffab;
mem[603]  = 80'h0010ffabffabffabffab;
mem[604]  = 80'h0010ffabffabffabffab;
mem[605]  = 80'h0010ffabffabffabffab;
mem[606]  = 80'h0010ffabffabffabffab;
mem[607]  = 80'h0010ffabffabffabffab;
mem[608]  = 80'h0010ffabffabffabffab;
mem[609]  = 80'h0010ffabffabffabffab;
mem[610]  = 80'h0010ffabffabffabffab;
mem[611]  = 80'h0010ffabffabffabffab;
mem[612]  = 80'h0010ffabffabffabffab;
mem[613]  = 80'h0010ffabffabffabffab;
mem[614]  = 80'h0010ffabffabffabffab;
mem[615]  = 80'h0010ffabffabffabffab;
mem[616]  = 80'h0010ffabffabffabffab;
mem[617]  = 80'h0010ffabffabffabffab;
mem[618]  = 80'h0010ffabffabffabffab;
mem[619]  = 80'h0010ffabffabffabffab;
mem[620]  = 80'h0010ffabffabffabffab;
mem[621]  = 80'h0010ffabffabffabffab;
mem[622]  = 80'h0010ffabffabffabffab;
mem[623]  = 80'h0010ffabffabffabffab;
mem[624]  = 80'h0010ffabffabffabffab;
mem[625]  = 80'h0010ffabffabffabffab;
mem[626]  = 80'h0010ffabffabffabffab;
mem[627]  = 80'h0010ffabffabffabffab;
mem[628]  = 80'h0010ffabffabffabffab;
mem[629]  = 80'h0010ffabffabffabffab;
mem[630]  = 80'h0010ffabffabffabffab;
mem[631]  = 80'h0010ffabffabffabffab;
mem[632]  = 80'h0010ffabffabffabffab;
mem[633]  = 80'h0010ffabffabffabffab;
mem[634]  = 80'h0010ffabffabffabffab;
mem[635]  = 80'h0010ffabffabffabffab;
mem[636]  = 80'h0010ffabffabffabffab;
mem[637]  = 80'h0010ffabffabffabffab;
mem[638]  = 80'h0010ffabffabffabffab;
mem[639]  = 80'h0010ffabffabffabffab;
mem[640]  = 80'h0010ffabffabffabffab;
mem[641]  = 80'h0010ffabffabffabffab;
mem[642]  = 80'h0010ffabffabffabffab;
mem[643]  = 80'h0010ffabffabffabffab;
mem[644]  = 80'h0010ffabffabffabffab;
mem[645]  = 80'h0010ffabffabffabffab;
mem[646]  = 80'h0010ffabffabffabffab;
mem[647]  = 80'h0010ffabffabffabffab;
mem[648]  = 80'h0010ffabffabffabffab;
mem[649]  = 80'h0010ffabffabffabffab;
mem[650]  = 80'h0010ffabffabffabffab;
mem[651]  = 80'h0010ffabffabffabffab;
mem[652]  = 80'h0010ffabffabffabffab;
mem[653]  = 80'h0010ffabffabffabffab;
mem[654]  = 80'h0010ffabffabffabffab;
mem[655]  = 80'h0010ffabffabffabffab;
mem[656]  = 80'h0010ffabffabffabffab;
mem[657]  = 80'h0010ffabffabffabffab;
mem[658]  = 80'h0010ffabffabffabffab;
mem[659]  = 80'h0010ffabffabffabffab;
mem[660]  = 80'h0010ffabffabffabffab;
mem[661]  = 80'h0010ffabffabffabffab;
mem[662]  = 80'h0010ffabffabffabffab;
mem[663]  = 80'h0010ffabffabffabffab;
mem[664]  = 80'h0010ffabffabffabffab;
mem[665]  = 80'h0010ffabffabffabffab;
mem[666]  = 80'h0010ffabffabffabffab;
mem[667]  = 80'h0010ffabffabffabffab;
mem[668]  = 80'h0010ffabffabffabffab;
mem[669]  = 80'h0010ffabffabffabffab;
mem[670]  = 80'h0010ffabffabffabffab;
mem[671]  = 80'h0010ffabffabffabffab;
mem[672]  = 80'h0010ffabffabffabffab;
mem[673]  = 80'h0010ffabffabffabffab;
mem[674]  = 80'h0010ffabffabffabffab;
mem[675]  = 80'h0010ffabffabffabffab;
mem[676]  = 80'h0010ffabffabffabffab;
mem[677]  = 80'h0010ffabffabffabffab;
mem[678]  = 80'h0010ffab61e70bff2fc3;
mem[679]  = 80'h001093c1a0c80b835d9d;
mem[680]  = 80'h0010d13ba6aa4cc505ba;
mem[681]  = 80'h0112cf5a000000000000;
mem[682]  = 80'h10100000010000010010;
mem[683]  = 80'h00109400000208004500;
mem[684]  = 80'h0010017f899f0000fffd;
mem[685]  = 80'h0010ae89c0550102c000;
mem[686]  = 80'h00100001ffabffabffab;
mem[687]  = 80'h0010ffabffabffabffab;
mem[688]  = 80'h0010ffabffabffabffab;
mem[689]  = 80'h0010ffabffabffabffab;
mem[690]  = 80'h0010ffabffabffabffab;
mem[691]  = 80'h0010ffabffabffabffab;
mem[692]  = 80'h0010ffabffabffabffab;
mem[693]  = 80'h0010ffabffabffabffab;
mem[694]  = 80'h0010ffabffabffabffab;
mem[695]  = 80'h0010ffabffabffabffab;
mem[696]  = 80'h0010ffabffabffabffab;
mem[697]  = 80'h0010ffabffabffabffab;
mem[698]  = 80'h0010ffabffabffabffab;
mem[699]  = 80'h0010ffabffabffabffab;
mem[700]  = 80'h0010ffabffabffabffab;
mem[701]  = 80'h0010ffabffabffabffab;
mem[702]  = 80'h0010ffabffabffabffab;
mem[703]  = 80'h0010ffabffabffabffab;
mem[704]  = 80'h0010ffabffabffabffab;
mem[705]  = 80'h0010ffabffabffabffab;
mem[706]  = 80'h0010ffabffabffabffab;
mem[707]  = 80'h0010ffabffabffabffab;
mem[708]  = 80'h0010ffabffabffabffab;
mem[709]  = 80'h0010ffabffabffabffab;
mem[710]  = 80'h0010ffabffabffabffab;
mem[711]  = 80'h0010ffabffabffabffab;
mem[712]  = 80'h0010ffabffabffabffab;
mem[713]  = 80'h0010ffabffabffabffab;
mem[714]  = 80'h0010ffabffabffabffab;
mem[715]  = 80'h0010ffabffabffabffab;
mem[716]  = 80'h0010ffabffabffabffab;
mem[717]  = 80'h0010ffabffabffabffab;
mem[718]  = 80'h0010ffabffabffabffab;
mem[719]  = 80'h0010ffabffabffabffab;
mem[720]  = 80'h0010ffabffabffabffab;
mem[721]  = 80'h0010ffabffabffabffab;
mem[722]  = 80'h0010ffabffabffabffab;
mem[723]  = 80'h0010ffabffabffabffab;
mem[724]  = 80'h0010ffabffabffabffab;
mem[725]  = 80'h0010ffabffabffabffab;
mem[726]  = 80'h0010ffabffabffabffab;
mem[727]  = 80'h0010ffabffabffabffab;
mem[728]  = 80'h0010ffabffabffabffab;
mem[729]  = 80'h0010ff6096d5d3f7ba51;
mem[730]  = 80'h00107e6b1a8c6ea87243;
mem[731]  = 80'h00106a407d5c7951ca29;
mem[732]  = 80'h01118800000000000000;
mem[733]  = 80'h10100000010000010010;
mem[734]  = 80'h00109400000208004500;
mem[735]  = 80'h001000d889a00000fffd;
mem[736]  = 80'h0010af2fc0550102c000;
mem[737]  = 80'h00100001ffabffabffab;
mem[738]  = 80'h0010ffabffabffabffab;
mem[739]  = 80'h0010ffabffabffabffab;
mem[740]  = 80'h0010ffabffabffabffab;
mem[741]  = 80'h0010ffabffabffabffab;
mem[742]  = 80'h0010ffabffabffabffab;
mem[743]  = 80'h0010ffabffabffabffab;
mem[744]  = 80'h0010ffabffabffabffab;
mem[745]  = 80'h0010ffabffabffabffab;
mem[746]  = 80'h0010ffabffabffabffab;
mem[747]  = 80'h0010ffabffabffabffab;
mem[748]  = 80'h0010ffabffabffabffab;
mem[749]  = 80'h0010ffabffabffabffab;
mem[750]  = 80'h0010ffabffabffabffab;
mem[751]  = 80'h0010ffabffabffabffab;
mem[752]  = 80'h0010ffabffabffabffab;
mem[753]  = 80'h0010ffabffabffabffab;
mem[754]  = 80'h0010ffabffabffabffab;
mem[755]  = 80'h0010ffabffabffabffab;
mem[756]  = 80'h0010ffabffabffabffab;
mem[757]  = 80'h0010ffabffabffabffab;
mem[758]  = 80'h0010ffabffabffabffab;
mem[759]  = 80'h0010ffab5fe5e8437673;
mem[760]  = 80'h00106044df5f908e8648;
mem[761]  = 80'h0010fef1e38308728fe0;
mem[762]  = 80'h01121bc1000000000000;
mem[763]  = 80'h10100000010000010010;
mem[764]  = 80'h00109400000208004500;
mem[765]  = 80'h0010035989a10000fffd;
mem[766]  = 80'h0010acadc0550102c000;
mem[767]  = 80'h00100001ffabffabffab;
mem[768]  = 80'h0010ffabffabffabffab;
mem[769]  = 80'h0010ffabffabffabffab;
mem[770]  = 80'h0010ffabffabffabffab;
mem[771]  = 80'h0010ffabffabffabffab;
mem[772]  = 80'h0010ffabffabffabffab;
mem[773]  = 80'h0010ffabffabffabffab;
mem[774]  = 80'h0010ffabffabffabffab;
mem[775]  = 80'h0010ffabffabffabffab;
mem[776]  = 80'h0010ffabffabffabffab;
mem[777]  = 80'h0010ffabffabffabffab;
mem[778]  = 80'h0010ffabffabffabffab;
mem[779]  = 80'h0010ffabffabffabffab;
mem[780]  = 80'h0010ffabffabffabffab;
mem[781]  = 80'h0010ffabffabffabffab;
mem[782]  = 80'h0010ffabffabffabffab;
mem[783]  = 80'h0010ffabffabffabffab;
mem[784]  = 80'h0010ffabffabffabffab;
mem[785]  = 80'h0010ffabffabffabffab;
mem[786]  = 80'h0010ffabffabffabffab;
mem[787]  = 80'h0010ffabffabffabffab;
mem[788]  = 80'h0010ffabffabffabffab;
mem[789]  = 80'h0010ffabffabffabffab;
mem[790]  = 80'h0010ffabffabffabffab;
mem[791]  = 80'h0010ffabffabffabffab;
mem[792]  = 80'h0010ffabffabffabffab;
mem[793]  = 80'h0010ffabffabffabffab;
mem[794]  = 80'h0010ffabffabffabffab;
mem[795]  = 80'h0010ffabffabffabffab;
mem[796]  = 80'h0010ffabffabffabffab;
mem[797]  = 80'h0010ffabffabffabffab;
mem[798]  = 80'h0010ffabffabffabffab;
mem[799]  = 80'h0010ffabffabffabffab;
mem[800]  = 80'h0010ffabffabffabffab;
mem[801]  = 80'h0010ffabffabffabffab;
mem[802]  = 80'h0010ffabffabffabffab;
mem[803]  = 80'h0010ffabffabffabffab;
mem[804]  = 80'h0010ffabffabffabffab;
mem[805]  = 80'h0010ffabffabffabffab;
mem[806]  = 80'h0010ffabffabffabffab;
mem[807]  = 80'h0010ffabffabffabffab;
mem[808]  = 80'h0010ffabffabffabffab;
mem[809]  = 80'h0010ffabffabffabffab;
mem[810]  = 80'h0010ffabffabffabffab;
mem[811]  = 80'h0010ffabffabffabffab;
mem[812]  = 80'h0010ffabffabffabffab;
mem[813]  = 80'h0010ffabffabffabffab;
mem[814]  = 80'h0010ffabffabffabffab;
mem[815]  = 80'h0010ffabffabffabffab;
mem[816]  = 80'h0010ffabffabffabffab;
mem[817]  = 80'h0010ffabffabffabffab;
mem[818]  = 80'h0010ffabffabffabffab;
mem[819]  = 80'h0010ffabffabffabffab;
mem[820]  = 80'h0010ffabffabffabffab;
mem[821]  = 80'h0010ffabffabffabffab;
mem[822]  = 80'h0010ffabffabffabffab;
mem[823]  = 80'h0010ffabffabffabffab;
mem[824]  = 80'h0010ffabffabffabffab;
mem[825]  = 80'h0010ffabffabffabffab;
mem[826]  = 80'h0010ffabffabffabffab;
mem[827]  = 80'h0010ffabffabffabffab;
mem[828]  = 80'h0010ffabffabffabffab;
mem[829]  = 80'h0010ffabffabffabffab;
mem[830]  = 80'h0010ffabffabffabffab;
mem[831]  = 80'h0010ffabffabffabffab;
mem[832]  = 80'h0010ffabffabffabffab;
mem[833]  = 80'h0010ffabffabffabffab;
mem[834]  = 80'h0010ffabffabffabffab;
mem[835]  = 80'h0010ffabffabffabffab;
mem[836]  = 80'h0010ffabffabffabffab;
mem[837]  = 80'h0010ffabffabffabffab;
mem[838]  = 80'h0010ffabffabffabffab;
mem[839]  = 80'h0010ffabffabffabffab;
mem[840]  = 80'h0010ffabffabffabffab;
mem[841]  = 80'h0010ffabffabffabffab;
mem[842]  = 80'h0010ffabffabffabffab;
mem[843]  = 80'h0010ffabffabffabffab;
mem[844]  = 80'h0010ffabffabffabffab;
mem[845]  = 80'h0010ffabffabffabffab;
mem[846]  = 80'h0010ffabffabffabffab;
mem[847]  = 80'h0010ffabffabffabffab;
mem[848]  = 80'h0010ffabffabffabffab;
mem[849]  = 80'h0010ffabffabffabffab;
mem[850]  = 80'h0010ffabffabffabffab;
mem[851]  = 80'h0010ffabffabffabffab;
mem[852]  = 80'h0010ffabffabffabffab;
mem[853]  = 80'h0010ffabffabffabffab;
mem[854]  = 80'h0010ffabffabffabffab;
mem[855]  = 80'h0010ffabffabffabffab;
mem[856]  = 80'h0010ffabffabffabffab;
mem[857]  = 80'h0010ffabffabffabffab;
mem[858]  = 80'h0010ffabffabffabffab;
mem[859]  = 80'h0010ffabffabffabffab;
mem[860]  = 80'h0010ffabffabffabffab;
mem[861]  = 80'h0010ffabffabffabffab;
mem[862]  = 80'h0010ffabffabffabffab;
mem[863]  = 80'h0010ffabffabffabffab;
mem[864]  = 80'h0010ffabffabffabffab;
mem[865]  = 80'h0010ffabffabffabffab;
mem[866]  = 80'h0010ffabffabffabffab;
mem[867]  = 80'h0010ffabffabffabffab;
mem[868]  = 80'h0010ffabffabffabffab;
mem[869]  = 80'h0010ffabff5e94366fae;
mem[870]  = 80'h00100aa2fb148d176373;
mem[871]  = 80'h001098c9a00e4ba281a5;
mem[872]  = 80'h01131bbb7d0000000000;
mem[873]  = 80'h10100000010000010010;
mem[874]  = 80'h00109400000208004500;
mem[875]  = 80'h001001c289a20000fffd;
mem[876]  = 80'h0010ae43c0550102c000;
mem[877]  = 80'h00100001ffabffabffab;
mem[878]  = 80'h0010ffabffabffabffab;
mem[879]  = 80'h0010ffabffabffabffab;
mem[880]  = 80'h0010ffabffabffabffab;
mem[881]  = 80'h0010ffabffabffabffab;
mem[882]  = 80'h0010ffabffabffabffab;
mem[883]  = 80'h0010ffabffabffabffab;
mem[884]  = 80'h0010ffabffabffabffab;
mem[885]  = 80'h0010ffabffabffabffab;
mem[886]  = 80'h0010ffabffabffabffab;
mem[887]  = 80'h0010ffabffabffabffab;
mem[888]  = 80'h0010ffabffabffabffab;
mem[889]  = 80'h0010ffabffabffabffab;
mem[890]  = 80'h0010ffabffabffabffab;
mem[891]  = 80'h0010ffabffabffabffab;
mem[892]  = 80'h0010ffabffabffabffab;
mem[893]  = 80'h0010ffabffabffabffab;
mem[894]  = 80'h0010ffabffabffabffab;
mem[895]  = 80'h0010ffabffabffabffab;
mem[896]  = 80'h0010ffabffabffabffab;
mem[897]  = 80'h0010ffabffabffabffab;
mem[898]  = 80'h0010ffabffabffabffab;
mem[899]  = 80'h0010ffabffabffabffab;
mem[900]  = 80'h0010ffabffabffabffab;
mem[901]  = 80'h0010ffabffabffabffab;
mem[902]  = 80'h0010ffabffabffabffab;
mem[903]  = 80'h0010ffabffabffabffab;
mem[904]  = 80'h0010ffabffabffabffab;
mem[905]  = 80'h0010ffabffabffabffab;
mem[906]  = 80'h0010ffabffabffabffab;
mem[907]  = 80'h0010ffabffabffabffab;
mem[908]  = 80'h0010ffabffabffabffab;
mem[909]  = 80'h0010ffabffabffabffab;
mem[910]  = 80'h0010ffabffabffabffab;
mem[911]  = 80'h0010ffabffabffabffab;
mem[912]  = 80'h0010ffabffabffabffab;
mem[913]  = 80'h0010ffabffabffabffab;
mem[914]  = 80'h0010ffabffabffabffab;
mem[915]  = 80'h0010ffabffabffabffab;
mem[916]  = 80'h0010ffabffabffabffab;
mem[917]  = 80'h0010ffabffabffabffab;
mem[918]  = 80'h0010ffabffabffabffab;
mem[919]  = 80'h0010ffabffabffabffab;
mem[920]  = 80'h0010ffabffabffabffab;
mem[921]  = 80'h0010ffabffabffabffab;
mem[922]  = 80'h0010ffabffabffabffab;
mem[923]  = 80'h0010ffabffabffabffab;
mem[924]  = 80'h0010ffabffabffabffab;
mem[925]  = 80'h0010ffabffabffabffab;
mem[926]  = 80'h0010ffabffabffabffab;
mem[927]  = 80'h0010ffabffabffabffab;
mem[928]  = 80'h0010ffabffab5d06541a;
mem[929]  = 80'h0010c680e53b48fa9f55;
mem[930]  = 80'h00106deb4452b8a04ff4;
mem[931]  = 80'h0114b4a5caac00000000;
mem[932]  = 80'h10100000010000010010;
mem[933]  = 80'h00109400000208004500;
mem[934]  = 80'h001003d189a30000fffd;
mem[935]  = 80'h0010ac33c0550102c000;
mem[936]  = 80'h00100001ffabffabffab;
mem[937]  = 80'h0010ffabffabffabffab;
mem[938]  = 80'h0010ffabffabffabffab;
mem[939]  = 80'h0010ffabffabffabffab;
mem[940]  = 80'h0010ffabffabffabffab;
mem[941]  = 80'h0010ffabffabffabffab;
mem[942]  = 80'h0010ffabffabffabffab;
mem[943]  = 80'h0010ffabffabffabffab;
mem[944]  = 80'h0010ffabffabffabffab;
mem[945]  = 80'h0010ffabffabffabffab;
mem[946]  = 80'h0010ffabffabffabffab;
mem[947]  = 80'h0010ffabffabffabffab;
mem[948]  = 80'h0010ffabffabffabffab;
mem[949]  = 80'h0010ffabffabffabffab;
mem[950]  = 80'h0010ffabffabffabffab;
mem[951]  = 80'h0010ffabffabffabffab;
mem[952]  = 80'h0010ffabffabffabffab;
mem[953]  = 80'h0010ffabffabffabffab;
mem[954]  = 80'h0010ffabffabffabffab;
mem[955]  = 80'h0010ffabffabffabffab;
mem[956]  = 80'h0010ffabffabffabffab;
mem[957]  = 80'h0010ffabffabffabffab;
mem[958]  = 80'h0010ffabffabffabffab;
mem[959]  = 80'h0010ffabffabffabffab;
mem[960]  = 80'h0010ffabffabffabffab;
mem[961]  = 80'h0010ffabffabffabffab;
mem[962]  = 80'h0010ffabffabffabffab;
mem[963]  = 80'h0010ffabffabffabffab;
mem[964]  = 80'h0010ffabffabffabffab;
mem[965]  = 80'h0010ffabffabffabffab;
mem[966]  = 80'h0010ffabffabffabffab;
mem[967]  = 80'h0010ffabffabffabffab;
mem[968]  = 80'h0010ffabffabffabffab;
mem[969]  = 80'h0010ffabffabffabffab;
mem[970]  = 80'h0010ffabffabffabffab;
mem[971]  = 80'h0010ffabffabffabffab;
mem[972]  = 80'h0010ffabffabffabffab;
mem[973]  = 80'h0010ffabffabffabffab;
mem[974]  = 80'h0010ffabffabffabffab;
mem[975]  = 80'h0010ffabffabffabffab;
mem[976]  = 80'h0010ffabffabffabffab;
mem[977]  = 80'h0010ffabffabffabffab;
mem[978]  = 80'h0010ffabffabffabffab;
mem[979]  = 80'h0010ffabffabffabffab;
mem[980]  = 80'h0010ffabffabffabffab;
mem[981]  = 80'h0010ffabffabffabffab;
mem[982]  = 80'h0010ffabffabffabffab;
mem[983]  = 80'h0010ffabffabffabffab;
mem[984]  = 80'h0010ffabffabffabffab;
mem[985]  = 80'h0010ffabffabffabffab;
mem[986]  = 80'h0010ffabffabffabffab;
mem[987]  = 80'h0010ffabffabffabffab;
mem[988]  = 80'h0010ffabffabffabffab;
mem[989]  = 80'h0010ffabffabffabffab;
mem[990]  = 80'h0010ffabffabffabffab;
mem[991]  = 80'h0010ffabffabffabffab;
mem[992]  = 80'h0010ffabffabffabffab;
mem[993]  = 80'h0010ffabffabffabffab;
mem[994]  = 80'h0010ffabffabffabffab;
mem[995]  = 80'h0010ffabffabffabffab;
mem[996]  = 80'h0010ffabffabffabffab;
mem[997]  = 80'h0010ffabffabffabffab;
mem[998]  = 80'h0010ffabffabffabffab;
mem[999]  = 80'h0010ffabffabffabffab;
mem[1000] = 80'h0010ffabffabffabffab;
mem[1001] = 80'h0010ffabffabffabffab;
mem[1002] = 80'h0010ffabffabffabffab;
mem[1003] = 80'h0010ffabffabffabffab;
mem[1004] = 80'h0010ffabffabffabffab;
mem[1005] = 80'h0010ffabffabffabffab;
mem[1006] = 80'h0010ffabffabffabffab;
mem[1007] = 80'h0010ffabffabffabffab;
mem[1008] = 80'h0010ffabffabffabffab;
mem[1009] = 80'h0010ffabffabffabffab;
mem[1010] = 80'h0010ffabffabffabffab;
mem[1011] = 80'h0010ffabffabffabffab;
mem[1012] = 80'h0010ffabffabffabffab;
mem[1013] = 80'h0010ffabffabffabffab;
mem[1014] = 80'h0010ffabffabffabffab;
mem[1015] = 80'h0010ffabffabffabffab;
mem[1016] = 80'h0010ffabffabffabffab;
mem[1017] = 80'h0010ffabffabffabffab;
mem[1018] = 80'h0010ffabffabffabffab;
mem[1019] = 80'h0010ffabffabffabffab;
mem[1020] = 80'h0010ffabffabffabffab;
mem[1021] = 80'h0010ffabffabffabffab;
mem[1022] = 80'h0010ffabffabffabffab;
mem[1023] = 80'h0010ffabffabffabffab;
mem[1024] = 80'h0010ffabffabffabffab;
mem[1025] = 80'h0010ffabffabffabffab;
mem[1026] = 80'h0010ffabffabffabffab;
mem[1027] = 80'h0010ffabffabffabffab;
mem[1028] = 80'h0010ffabffabffabffab;
mem[1029] = 80'h0010ffabffabffabffab;
mem[1030] = 80'h0010ffabffabffabffab;
mem[1031] = 80'h0010ffabffabffabffab;
mem[1032] = 80'h0010ffabffabffabffab;
mem[1033] = 80'h0010ffabffabffabffab;
mem[1034] = 80'h0010ffabffabffabffab;
mem[1035] = 80'h0010ffabffabffabffab;
mem[1036] = 80'h0010ffabffabffabffab;
mem[1037] = 80'h0010ffabffabffabffab;
mem[1038] = 80'h0010ffabffabffabffab;
mem[1039] = 80'h0010ffabffabffabffab;
mem[1040] = 80'h0010ffabffabffabffab;
mem[1041] = 80'h0010ffabffabffabffab;
mem[1042] = 80'h0010ffabffabffabffab;
mem[1043] = 80'h0010ffabffabffabffab;
mem[1044] = 80'h0010ffabffabffabffab;
mem[1045] = 80'h0010ffabffabffabffab;
mem[1046] = 80'h0010ffabffabffabffab;
mem[1047] = 80'h0010ffabffabffabffab;
mem[1048] = 80'h0010ffabffabffabffab;
mem[1049] = 80'h0010ffabffabffabffab;
mem[1050] = 80'h0010ffabffabffabffab;
mem[1051] = 80'h0010ffabffabffabffab;
mem[1052] = 80'h0010ffabffabffabffab;
mem[1053] = 80'h0010ffabff5c778a361e;
mem[1054] = 80'h0010f92784832818b898;
mem[1055] = 80'h00103a4003329e2c1818;
mem[1056] = 80'h011315868d0000000000;
mem[1057] = 80'h10100000010000010010;
mem[1058] = 80'h00109400000208004500;
mem[1059] = 80'h001001fe89a40000fffd;
mem[1060] = 80'h0010ae05c0550102c000;
mem[1061] = 80'h00100001ffabffabffab;
mem[1062] = 80'h0010ffabffabffabffab;
mem[1063] = 80'h0010ffabffabffabffab;
mem[1064] = 80'h0010ffabffabffabffab;
mem[1065] = 80'h0010ffabffabffabffab;
mem[1066] = 80'h0010ffabffabffabffab;
mem[1067] = 80'h0010ffabffabffabffab;
mem[1068] = 80'h0010ffabffabffabffab;
mem[1069] = 80'h0010ffabffabffabffab;
mem[1070] = 80'h0010ffabffabffabffab;
mem[1071] = 80'h0010ffabffabffabffab;
mem[1072] = 80'h0010ffabffabffabffab;
mem[1073] = 80'h0010ffabffabffabffab;
mem[1074] = 80'h0010ffabffabffabffab;
mem[1075] = 80'h0010ffabffabffabffab;
mem[1076] = 80'h0010ffabffabffabffab;
mem[1077] = 80'h0010ffabffabffabffab;
mem[1078] = 80'h0010ffabffabffabffab;
mem[1079] = 80'h0010ffabffabffabffab;
mem[1080] = 80'h0010ffabffabffabffab;
mem[1081] = 80'h0010ffabffabffabffab;
mem[1082] = 80'h0010ffabffabffabffab;
mem[1083] = 80'h0010ffabffabffabffab;
mem[1084] = 80'h0010ffabffabffabffab;
mem[1085] = 80'h0010ffabffabffabffab;
mem[1086] = 80'h0010ffabffabffabffab;
mem[1087] = 80'h0010ffabffabffabffab;
mem[1088] = 80'h0010ffabffabffabffab;
mem[1089] = 80'h0010ffabffabffabffab;
mem[1090] = 80'h0010ffabffabffabffab;
mem[1091] = 80'h0010ffabffabffabffab;
mem[1092] = 80'h0010ffabffabffabffab;
mem[1093] = 80'h0010ffabffabffabffab;
mem[1094] = 80'h0010ffabffabffabffab;
mem[1095] = 80'h0010ffabffabffabffab;
mem[1096] = 80'h0010ffabffabffabffab;
mem[1097] = 80'h0010ffabffabffabffab;
mem[1098] = 80'h0010ffabffabffabffab;
mem[1099] = 80'h0010ffabffabffabffab;
mem[1100] = 80'h0010ffabffabffabffab;
mem[1101] = 80'h0010ffabffabffabffab;
mem[1102] = 80'h0010ffabffabffabffab;
mem[1103] = 80'h0010ffabffabffabffab;
mem[1104] = 80'h0010ffabffabffabffab;
mem[1105] = 80'h0010ffabffabffabffab;
mem[1106] = 80'h0010ffabffabffabffab;
mem[1107] = 80'h0010ffabffabffabffab;
mem[1108] = 80'h0010ffabffabffabffab;
mem[1109] = 80'h0010ffabffabffabffab;
mem[1110] = 80'h0010ffabffabffabffab;
mem[1111] = 80'h0010ffabffabffabffab;
mem[1112] = 80'h0010ffabffabffabffab;
mem[1113] = 80'h0010ffabffabffabffab;
mem[1114] = 80'h0010ffabffabffabffab;
mem[1115] = 80'h0010ffabffabffabffab;
mem[1116] = 80'h0010ffabffabffabffab;
mem[1117] = 80'h0010ffabffabffabffab;
mem[1118] = 80'h0010ffabffabffabffab;
mem[1119] = 80'h0010ffabffabffabffab;
mem[1120] = 80'h00105b534edccfeda804;
mem[1121] = 80'h00103bc709d4a4dc52e6;
mem[1122] = 80'h01109740093fc006df3e;
mem[1123] = 80'h10100000010000010010;
mem[1124] = 80'h00109400000208004500;
mem[1125] = 80'h0010011689a50000fffd;
mem[1126] = 80'h0010aeecc0550102c000;
mem[1127] = 80'h00100001ffabffabffab;
mem[1128] = 80'h0010ffabffabffabffab;
mem[1129] = 80'h0010ffabffabffabffab;
mem[1130] = 80'h0010ffabffabffabffab;
mem[1131] = 80'h0010ffabffabffabffab;
mem[1132] = 80'h0010ffabffabffabffab;
mem[1133] = 80'h0010ffabffabffabffab;
mem[1134] = 80'h0010ffabffabffabffab;
mem[1135] = 80'h0010ffabffabffabffab;
mem[1136] = 80'h0010ffabffabffabffab;
mem[1137] = 80'h0010ffabffabffabffab;
mem[1138] = 80'h0010ffabffabffabffab;
mem[1139] = 80'h0010ffabffabffabffab;
mem[1140] = 80'h0010ffabffabffabffab;
mem[1141] = 80'h0010ffabffabffabffab;
mem[1142] = 80'h0010ffabffabffabffab;
mem[1143] = 80'h0010ffabffabffabffab;
mem[1144] = 80'h0010ffabffabffabffab;
mem[1145] = 80'h0010ffabffabffabffab;
mem[1146] = 80'h0010ffabffabffabffab;
mem[1147] = 80'h0010ffabffabffabffab;
mem[1148] = 80'h0010ffabffabffabffab;
mem[1149] = 80'h0010ffabffabffabffab;
mem[1150] = 80'h0010ffabffabffabffab;
mem[1151] = 80'h0010ffabffabffabffab;
mem[1152] = 80'h0010ffabffabffabffab;
mem[1153] = 80'h0010ffabffabffabffab;
mem[1154] = 80'h0010ffabffabffabffab;
mem[1155] = 80'h0010ffabffabffabffab;
mem[1156] = 80'h0010ffabffabffabffab;
mem[1157] = 80'h00105a2290f017946abb;
mem[1158] = 80'h0010f0158e39510d67b7;
mem[1159] = 80'h01102bda2fafd3b4178b;
mem[1160] = 80'h10100000010000010010;
mem[1161] = 80'h00109400000208004500;
mem[1162] = 80'h001000a289a60000fffd;
mem[1163] = 80'h0010af5fc0550102c000;
mem[1164] = 80'h00100001ffabffabffab;
mem[1165] = 80'h0010ffabffabffabffab;
mem[1166] = 80'h0010ffabffabffabffab;
mem[1167] = 80'h0010ffabffabffabffab;
mem[1168] = 80'h0010ffabffabffabffab;
mem[1169] = 80'h0010ffabffabffabffab;
mem[1170] = 80'h0010ffabffabffabffab;
mem[1171] = 80'h0010ffabffabffabffab;
mem[1172] = 80'h0010ffabffabffabffab;
mem[1173] = 80'h0010ffabffabffabffab;
mem[1174] = 80'h0010ffabffabffabffab;
mem[1175] = 80'h0010ffabffabffabffab;
mem[1176] = 80'h0010ffabffabffabffab;
mem[1177] = 80'h0010ffabffabffabffab;
mem[1178] = 80'h0010ffabffabffabffab;
mem[1179] = 80'h0010ffabffab59b0f285;
mem[1180] = 80'h00107f1e2d7bac62060f;
mem[1181] = 80'h00104f7daf4536581fa3;
mem[1182] = 80'h0114acf0ac8c00000000;
mem[1183] = 80'h10100000010000010010;
mem[1184] = 80'h00109400000208004500;
mem[1185] = 80'h0010006989a70000fffd;
mem[1186] = 80'h0010af97c0550102c000;
mem[1187] = 80'h00100001ffabffabffab;
mem[1188] = 80'h0010ffabffabffabffab;
mem[1189] = 80'h0010ffabffabffabffab;
mem[1190] = 80'h0010ffabffabffabffab;
mem[1191] = 80'h0010ffabffabffabffab;
mem[1192] = 80'h0010ffabffabffabffab;
mem[1193] = 80'h0010ffabffabffabffab;
mem[1194] = 80'h0010ffabffabffabffab;
mem[1195] = 80'h0010ffabff58c12ca9a7;
mem[1196] = 80'h001067efc467b081e2ba;
mem[1197] = 80'h0010ad14148565a5ae6f;
mem[1198] = 80'h0113a818640000000000;
mem[1199] = 80'h10100000010000010010;
mem[1200] = 80'h00109400000208004500;
mem[1201] = 80'h0010032489a80000fffd;
mem[1202] = 80'h0010acdbc0550102c000;
mem[1203] = 80'h00100001ffabffabffab;
mem[1204] = 80'h0010ffabffabffabffab;
mem[1205] = 80'h0010ffabffabffabffab;
mem[1206] = 80'h0010ffabffabffabffab;
mem[1207] = 80'h0010ffabffabffabffab;
mem[1208] = 80'h0010ffabffabffabffab;
mem[1209] = 80'h0010ffabffabffabffab;
mem[1210] = 80'h0010ffabffabffabffab;
mem[1211] = 80'h0010ffabffabffabffab;
mem[1212] = 80'h0010ffabffabffabffab;
mem[1213] = 80'h0010ffabffabffabffab;
mem[1214] = 80'h0010ffabffabffabffab;
mem[1215] = 80'h0010ffabffabffabffab;
mem[1216] = 80'h0010ffabffabffabffab;
mem[1217] = 80'h0010ffabffabffabffab;
mem[1218] = 80'h0010ffabffabffabffab;
mem[1219] = 80'h0010ffabffabffabffab;
mem[1220] = 80'h0010ffabffabffabffab;
mem[1221] = 80'h0010ffabffabffabffab;
mem[1222] = 80'h0010ffabffabffabffab;
mem[1223] = 80'h0010ffabffabffabffab;
mem[1224] = 80'h0010ffabffabffabffab;
mem[1225] = 80'h0010ffabffabffabffab;
mem[1226] = 80'h0010ffabffabffabffab;
mem[1227] = 80'h0010ffabffabffabffab;
mem[1228] = 80'h0010ffabffabffabffab;
mem[1229] = 80'h0010ffabffabffabffab;
mem[1230] = 80'h0010ffabffabffabffab;
mem[1231] = 80'h0010ffabffabffabffab;
mem[1232] = 80'h0010ffabffabffabffab;
mem[1233] = 80'h0010ffabffabffabffab;
mem[1234] = 80'h0010ffabffabffabffab;
mem[1235] = 80'h0010ffabffabffabffab;
mem[1236] = 80'h0010ffabffabffabffab;
mem[1237] = 80'h0010ffabffabffabffab;
mem[1238] = 80'h0010ffabffabffabffab;
mem[1239] = 80'h0010ffabffabffabffab;
mem[1240] = 80'h0010ffabffabffabffab;
mem[1241] = 80'h0010ffabffabffabffab;
mem[1242] = 80'h0010ffabffabffabffab;
mem[1243] = 80'h0010ffabffabffabffab;
mem[1244] = 80'h0010ffabffabffabffab;
mem[1245] = 80'h0010ffabffabffabffab;
mem[1246] = 80'h0010ffabffabffabffab;
mem[1247] = 80'h0010ffabffabffabffab;
mem[1248] = 80'h0010ffabffabffabffab;
mem[1249] = 80'h0010ffabffabffabffab;
mem[1250] = 80'h0010ffabffabffabffab;
mem[1251] = 80'h0010ffabffabffabffab;
mem[1252] = 80'h0010ffabffabffabffab;
mem[1253] = 80'h0010ffabffabffabffab;
mem[1254] = 80'h0010ffabffabffabffab;
mem[1255] = 80'h0010ffabffabffabffab;
mem[1256] = 80'h0010ffabffabffabffab;
mem[1257] = 80'h0010ffabffabffabffab;
mem[1258] = 80'h0010ffabffabffabffab;
mem[1259] = 80'h0010ffabffabffabffab;
mem[1260] = 80'h0010ffabffabffabffab;
mem[1261] = 80'h0010ffabffabffabffab;
mem[1262] = 80'h0010ffabffabffabffab;
mem[1263] = 80'h0010ffabffabffabffab;
mem[1264] = 80'h0010ffabffabffabffab;
mem[1265] = 80'h0010ffabffabffabffab;
mem[1266] = 80'h0010ffabffabffabffab;
mem[1267] = 80'h0010ffabffabffabffab;
mem[1268] = 80'h0010ffabffabffabffab;
mem[1269] = 80'h0010ffabffabffabffab;
mem[1270] = 80'h0010ffabffabffabffab;
mem[1271] = 80'h0010ffabffabffabffab;
mem[1272] = 80'h0010ffabffabffabffab;
mem[1273] = 80'h0010ffabffabffabffab;
mem[1274] = 80'h0010ffabffabffabffab;
mem[1275] = 80'h0010ffabffabffabffab;
mem[1276] = 80'h0010ffabffabffabffab;
mem[1277] = 80'h0010ffabffabffabffab;
mem[1278] = 80'h0010ffabffabffabffab;
mem[1279] = 80'h0010ffabffabffabffab;
mem[1280] = 80'h0010ffabffabffabffab;
mem[1281] = 80'h0010ffabffabffabffab;
mem[1282] = 80'h0010ffabffabffabffab;
mem[1283] = 80'h0010ffabffabffabffab;
mem[1284] = 80'h0010ffabffabffabffab;
mem[1285] = 80'h0010ffabffabffabffab;
mem[1286] = 80'h0010ffabffabffabffab;
mem[1287] = 80'h0010ffabffabffabffab;
mem[1288] = 80'h0010ffabffabffabffab;
mem[1289] = 80'h0010ffabffabffabffab;
mem[1290] = 80'h0010ffabffabffabffab;
mem[1291] = 80'h0010ffabffabffabffab;
mem[1292] = 80'h0010ffabffabffabffab;
mem[1293] = 80'h0010ffabffabffabffab;
mem[1294] = 80'h0010ffabffabffabffab;
mem[1295] = 80'h0010ffabffabffabffab;
mem[1296] = 80'h0010ffabffabffabffab;
mem[1297] = 80'h0010ffabffabffabffab;
mem[1298] = 80'h0010ffabffabffab57f9;
mem[1299] = 80'h00107b50dd37327addbc;
mem[1300] = 80'h001024d736bfa08e8fc8;
mem[1301] = 80'h0116b359fc4c47a60000;
mem[1302] = 80'h10100000010000010010;
mem[1303] = 80'h00109400000208004500;
mem[1304] = 80'h0010048089a90000fffd;
mem[1305] = 80'h0010ab7ec0550102c000;
mem[1306] = 80'h00100001ffabffabffab;
mem[1307] = 80'h0010ffabffabffabffab;
mem[1308] = 80'h0010ffabffabffabffab;
mem[1309] = 80'h0010ffabffabffabffab;
mem[1310] = 80'h0010ffabffabffabffab;
mem[1311] = 80'h0010ffabffabffabffab;
mem[1312] = 80'h0010ffabffabffabffab;
mem[1313] = 80'h0010ffabffabffabffab;
mem[1314] = 80'h0010ffabffabffabffab;
mem[1315] = 80'h0010ffabffabffabffab;
mem[1316] = 80'h0010ffabffabffabffab;
mem[1317] = 80'h0010ffabffabffabffab;
mem[1318] = 80'h0010ffabffabffabffab;
mem[1319] = 80'h0010ffabffabffabffab;
mem[1320] = 80'h0010ffabffabffabffab;
mem[1321] = 80'h0010ffabffabffabffab;
mem[1322] = 80'h0010ffabffabffabffab;
mem[1323] = 80'h0010ffabffabffabffab;
mem[1324] = 80'h0010ffabffabffabffab;
mem[1325] = 80'h0010ffabffabffabffab;
mem[1326] = 80'h0010ffabffabffabffab;
mem[1327] = 80'h0010ffabffabffabffab;
mem[1328] = 80'h0010ffabffabffabffab;
mem[1329] = 80'h0010ffabffabffabffab;
mem[1330] = 80'h0010ffabffabffabffab;
mem[1331] = 80'h0010ffabffabffabffab;
mem[1332] = 80'h0010ffabffabffabffab;
mem[1333] = 80'h0010ffabffabffabffab;
mem[1334] = 80'h0010ffabffabffabffab;
mem[1335] = 80'h0010ffabffabffabffab;
mem[1336] = 80'h0010ffabffabffabffab;
mem[1337] = 80'h0010ffabffabffabffab;
mem[1338] = 80'h0010ffabffabffabffab;
mem[1339] = 80'h0010ffabffabffabffab;
mem[1340] = 80'h0010ffabffabffabffab;
mem[1341] = 80'h0010ffabffabffabffab;
mem[1342] = 80'h0010ffabffabffabffab;
mem[1343] = 80'h0010ffabffabffabffab;
mem[1344] = 80'h0010ffabffabffabffab;
mem[1345] = 80'h0010ffabffabffabffab;
mem[1346] = 80'h0010ffabffabffabffab;
mem[1347] = 80'h0010ffabffabffabffab;
mem[1348] = 80'h0010ffabffabffabffab;
mem[1349] = 80'h0010ffabffabffabffab;
mem[1350] = 80'h0010ffabffabffabffab;
mem[1351] = 80'h0010ffabffabffabffab;
mem[1352] = 80'h0010ffabffabffabffab;
mem[1353] = 80'h0010ffabffabffabffab;
mem[1354] = 80'h0010ffabffabffabffab;
mem[1355] = 80'h0010ffabffabffabffab;
mem[1356] = 80'h0010ffabffabffabffab;
mem[1357] = 80'h0010ffabffabffabffab;
mem[1358] = 80'h0010ffabffabffabffab;
mem[1359] = 80'h0010ffabffabffabffab;
mem[1360] = 80'h0010ffabffabffabffab;
mem[1361] = 80'h0010ffabffabffabffab;
mem[1362] = 80'h0010ffabffabffabffab;
mem[1363] = 80'h0010ffabffabffabffab;
mem[1364] = 80'h0010ffabffabffabffab;
mem[1365] = 80'h0010ffabffabffabffab;
mem[1366] = 80'h0010ffabffabffabffab;
mem[1367] = 80'h0010ffabffabffabffab;
mem[1368] = 80'h0010ffabffabffabffab;
mem[1369] = 80'h0010ffabffabffabffab;
mem[1370] = 80'h0010ffabffabffabffab;
mem[1371] = 80'h0010ffabffabffabffab;
mem[1372] = 80'h0010ffabffabffabffab;
mem[1373] = 80'h0010ffabffabffabffab;
mem[1374] = 80'h0010ffabffabffabffab;
mem[1375] = 80'h0010ffabffabffabffab;
mem[1376] = 80'h0010ffabffabffabffab;
mem[1377] = 80'h0010ffabffabffabffab;
mem[1378] = 80'h0010ffabffabffabffab;
mem[1379] = 80'h0010ffabffabffabffab;
mem[1380] = 80'h0010ffabffabffabffab;
mem[1381] = 80'h0010ffabffabffabffab;
mem[1382] = 80'h0010ffabffabffabffab;
mem[1383] = 80'h0010ffabffabffabffab;
mem[1384] = 80'h0010ffabffabffabffab;
mem[1385] = 80'h0010ffabffabffabffab;
mem[1386] = 80'h0010ffabffabffabffab;
mem[1387] = 80'h0010ffabffabffabffab;
mem[1388] = 80'h0010ffabffabffabffab;
mem[1389] = 80'h0010ffabffabffabffab;
mem[1390] = 80'h0010ffabffabffabffab;
mem[1391] = 80'h0010ffabffabffabffab;
mem[1392] = 80'h0010ffabffabffabffab;
mem[1393] = 80'h0010ffabffabffabffab;
mem[1394] = 80'h0010ffabffabffabffab;
mem[1395] = 80'h0010ffabffabffabffab;
mem[1396] = 80'h0010ffabffabffabffab;
mem[1397] = 80'h0010ffabffabffabffab;
mem[1398] = 80'h0010ffabffabffabffab;
mem[1399] = 80'h0010ffabffabffabffab;
mem[1400] = 80'h0010ffabffabffabffab;
mem[1401] = 80'h0010ffabffabffabffab;
mem[1402] = 80'h0010ffabffabffabffab;
mem[1403] = 80'h0010ffabffabffabffab;
mem[1404] = 80'h0010ffabffabffabffab;
mem[1405] = 80'h0010ffabffabffabffab;
mem[1406] = 80'h0010ffabffabffabffab;
mem[1407] = 80'h0010ffabffabffabffab;
mem[1408] = 80'h0010ffabffabffabffab;
mem[1409] = 80'h0010ffabffabffabffab;
mem[1410] = 80'h0010ffabffabffabffab;
mem[1411] = 80'h0010ffabffabffabffab;
mem[1412] = 80'h0010ffabffabffabffab;
mem[1413] = 80'h0010ffabffabffabffab;
mem[1414] = 80'h0010ffabffabffabffab;
mem[1415] = 80'h0010ffabffabffabffab;
mem[1416] = 80'h0010ffabffabffabffab;
mem[1417] = 80'h0010ffabffabffabffab;
mem[1418] = 80'h0010ffabffabffabffab;
mem[1419] = 80'h0010ffabffabffabffab;
mem[1420] = 80'h0010ffabffabffabffab;
mem[1421] = 80'h0010ffabffabffabffab;
mem[1422] = 80'h0010ffabffabffabffab;
mem[1423] = 80'h0010ffabffabffabffab;
mem[1424] = 80'h0010ffabffabffabffab;
mem[1425] = 80'h0010ffabffabffabffab;
mem[1426] = 80'h0010ffabffabffabffab;
mem[1427] = 80'h0010ffabffabffabffab;
mem[1428] = 80'h0010ffabffabffabffab;
mem[1429] = 80'h0010ffabffabffabffab;
mem[1430] = 80'h0010ffabffabffabffab;
mem[1431] = 80'h0010ffabffabffabffab;
mem[1432] = 80'h0010ffabffabffabffab;
mem[1433] = 80'h0010ffabffabffabffab;
mem[1434] = 80'h0010ffabffabffabffab;
mem[1435] = 80'h0010ffabffabffabffab;
mem[1436] = 80'h0010ffabffabffabffab;
mem[1437] = 80'h0010ffabffabffabffab;
mem[1438] = 80'h0010ffabffabffabffab;
mem[1439] = 80'h0010ffabffabffabffab;
mem[1440] = 80'h0010ffabffabffabffab;
mem[1441] = 80'h0010ffabffabffabffab;
mem[1442] = 80'h0010ffabffabffabffab;
mem[1443] = 80'h0010ffabffabffabffab;
mem[1444] = 80'h0010ffabffabffabffab;
mem[1445] = 80'h0010ffab5688a57c054e;
mem[1446] = 80'h0010f0c5166ea33ac36c;
mem[1447] = 80'h0010f0dfa9edf60373a0;
mem[1448] = 80'h0112ab8d000000000000;
mem[1449] = 80'h00000000000000000000;
mem[1450] = 80'h00000000000000000000;
mem[1451] = 80'h00000000000000000000;
mem[1452] = 80'h00000000000000000000;
mem[1453] = 80'h00000000000000000000;
mem[1454] = 80'h00000000000000000000;
mem[1455] = 80'h00000000000000000000;
mem[1456] = 80'h00000000000000000000;
mem[1457] = 80'h00000000000000000000;
mem[1458] = 80'h00000000000000000000;
mem[1459] = 80'h00000000000000000000;
mem[1460] = 80'h00000000000000000000;
mem[1461] = 80'h00000000000000000000;
mem[1462] = 80'h00000000000000000000;
mem[1463] = 80'h00000000000000000000;
mem[1464] = 80'h00000000000000000000;
mem[1465] = 80'h00000000000000000000;
mem[1466] = 80'h00000000000000000000;
mem[1467] = 80'h00000000000000000000;
mem[1468] = 80'h00000000000000000000;
mem[1469] = 80'h00000000000000000000;
mem[1470] = 80'h00000000000000000000;
mem[1471] = 80'h10100000010000010010;
mem[1472] = 80'h00109400000208004500;
mem[1473] = 80'h0010052e89aa0000fffd;
mem[1474] = 80'h0010aacfc0550102c000;
mem[1475] = 80'h00100001ffabffabffab;
mem[1476] = 80'h0010ffabffabffabffab;
mem[1477] = 80'h0010ffabffabffabffab;
mem[1478] = 80'h0010ffabffabffabffab;
mem[1479] = 80'h0010ffabffabffabffab;
mem[1480] = 80'h0010ffabffabffabffab;
mem[1481] = 80'h0010ffabffabffabffab;
mem[1482] = 80'h0010ffabffabffabffab;
mem[1483] = 80'h0010ffabffabffabffab;
mem[1484] = 80'h0010ffabffabffabffab;
mem[1485] = 80'h0010ffabffabffabffab;
mem[1486] = 80'h0010ffabffabffabffab;
mem[1487] = 80'h0010ffabffabffabffab;
mem[1488] = 80'h0010ffabffabffabffab;
mem[1489] = 80'h0010ffabffabffabffab;
mem[1490] = 80'h0010ffabffabffabffab;
mem[1491] = 80'h0010ffabffabffabffab;
mem[1492] = 80'h0010ffabffabffabffab;
mem[1493] = 80'h0010ffabffabffabffab;
mem[1494] = 80'h0010ffabffabffabffab;
mem[1495] = 80'h0010ffabffabffabffab;
mem[1496] = 80'h0010ffabffabffabffab;
mem[1497] = 80'h0010ffabffabffabffab;
mem[1498] = 80'h0010ffabffabffabffab;
mem[1499] = 80'h0010ffabffabffabffab;
mem[1500] = 80'h0010ffabffabffabffab;
mem[1501] = 80'h0010ffabffabffabffab;
mem[1502] = 80'h0010ffabffabffabffab;
mem[1503] = 80'h0010ffabffabffabffab;
mem[1504] = 80'h0010ffabffabffabffab;
mem[1505] = 80'h0010ffabffabffabffab;
mem[1506] = 80'h0010ffabffabffabffab;
mem[1507] = 80'h0010ffabffabffabffab;
mem[1508] = 80'h0010ffabffabffabffab;
mem[1509] = 80'h0010ffabffabffabffab;
mem[1510] = 80'h0010ffabffabffabffab;
mem[1511] = 80'h0010ffabffabffabffab;
mem[1512] = 80'h0010ffabffabffabffab;
mem[1513] = 80'h0010ffabffabffabffab;
mem[1514] = 80'h0010ffabffabffabffab;
mem[1515] = 80'h0010ffabffabffabffab;
mem[1516] = 80'h0010ffabffabffabffab;
mem[1517] = 80'h0010ffabffabffabffab;
mem[1518] = 80'h0010ffabffabffabffab;
mem[1519] = 80'h0010ffabffabffabffab;
mem[1520] = 80'h0010ffabffabffabffab;
mem[1521] = 80'h0010ffabffabffabffab;
mem[1522] = 80'h0010ffabffabffabffab;
mem[1523] = 80'h0010ffabffabffabffab;
mem[1524] = 80'h0010ffabffabffabffab;
mem[1525] = 80'h0010ffabffabffabffab;
mem[1526] = 80'h0010ffabffabffabffab;
mem[1527] = 80'h0010ffabffabffabffab;
mem[1528] = 80'h0010ffabffabffabffab;
mem[1529] = 80'h0010ffabffabffabffab;
mem[1530] = 80'h0010ffabffabffabffab;
mem[1531] = 80'h0010ffabffabffabffab;
mem[1532] = 80'h0010ffabffabffabffab;
mem[1533] = 80'h0010ffabffabffabffab;
mem[1534] = 80'h0010ffabffabffabffab;
mem[1535] = 80'h0010ffabffabffabffab;
mem[1536] = 80'h0010ffabffabffabffab;
mem[1537] = 80'h0010ffabffabffabffab;
mem[1538] = 80'h0010ffabffabffabffab;
mem[1539] = 80'h0010ffabffabffabffab;
mem[1540] = 80'h0010ffabffabffabffab;
mem[1541] = 80'h0010ffabffabffabffab;
mem[1542] = 80'h0010ffabffabffabffab;
mem[1543] = 80'h0010ffabffabffabffab;
mem[1544] = 80'h0010ffabffabffabffab;
mem[1545] = 80'h0010ffabffabffabffab;
mem[1546] = 80'h0010ffabffabffabffab;
mem[1547] = 80'h0010ffabffabffabffab;
mem[1548] = 80'h0010ffabffabffabffab;
mem[1549] = 80'h0010ffabffabffabffab;
mem[1550] = 80'h0010ffabffabffabffab;
mem[1551] = 80'h0010ffabffabffabffab;
mem[1552] = 80'h0010ffabffabffabffab;
mem[1553] = 80'h0010ffabffabffabffab;
mem[1554] = 80'h0010ffabffabffabffab;
mem[1555] = 80'h0010ffabffabffabffab;
mem[1556] = 80'h0010ffabffabffabffab;
mem[1557] = 80'h0010ffabffabffabffab;
mem[1558] = 80'h0010ffabffabffabffab;
mem[1559] = 80'h0010ffabffabffabffab;
mem[1560] = 80'h0010ffabffabffabffab;
mem[1561] = 80'h0010ffabffabffabffab;
mem[1562] = 80'h0010ffabffabffabffab;
mem[1563] = 80'h0010ffabffabffabffab;
mem[1564] = 80'h0010ffabffabffabffab;
mem[1565] = 80'h0010ffabffabffabffab;
mem[1566] = 80'h0010ffabffabffabffab;
mem[1567] = 80'h0010ffabffabffabffab;
mem[1568] = 80'h0010ffabffabffabffab;
mem[1569] = 80'h0010ffabffabffabffab;
mem[1570] = 80'h0010ffabffabffabffab;
mem[1571] = 80'h0010ffabffabffabffab;
mem[1572] = 80'h0010ffabffabffabffab;
mem[1573] = 80'h0010ffabffabffabffab;
mem[1574] = 80'h0010ffabffabffabffab;
mem[1575] = 80'h0010ffabffabffabffab;
mem[1576] = 80'h0010ffabffabffabffab;
mem[1577] = 80'h0010ffabffabffabffab;
mem[1578] = 80'h0010ffabffabffabffab;
mem[1579] = 80'h0010ffabffabffabffab;
mem[1580] = 80'h0010ffabffabffabffab;
mem[1581] = 80'h0010ffabffabffabffab;
mem[1582] = 80'h0010ffabffabffabffab;
mem[1583] = 80'h0010ffabffabffabffab;
mem[1584] = 80'h0010ffabffabffabffab;
mem[1585] = 80'h0010ffabffabffabffab;
mem[1586] = 80'h0010ffabffabffabffab;
mem[1587] = 80'h0010ffabffabffabffab;
mem[1588] = 80'h0010ffabffabffabffab;
mem[1589] = 80'h0010ffabffabffabffab;
mem[1590] = 80'h0010ffabffabffabffab;
mem[1591] = 80'h0010ffabffabffabffab;
mem[1592] = 80'h0010ffabffabffabffab;
mem[1593] = 80'h0010ffabffabffabffab;
mem[1594] = 80'h0010ffabffabffabffab;
mem[1595] = 80'h0010ffabffabffabffab;
mem[1596] = 80'h0010ffabffabffabffab;
mem[1597] = 80'h0010ffabffabffabffab;
mem[1598] = 80'h0010ffabffabffabffab;
mem[1599] = 80'h0010ffabffabffabffab;
mem[1600] = 80'h0010ffabffabffabffab;
mem[1601] = 80'h0010ffabffabffabffab;
mem[1602] = 80'h0010ffabffabffabffab;
mem[1603] = 80'h0010ffabffabffabffab;
mem[1604] = 80'h0010ffabffabffabffab;
mem[1605] = 80'h0010ffabffabffabffab;
mem[1606] = 80'h0010ffabffabffabffab;
mem[1607] = 80'h0010ffabffabffabffab;
mem[1608] = 80'h0010ffabffabffabffab;
mem[1609] = 80'h0010ffabffabffabffab;
mem[1610] = 80'h0010ffabffabffabffab;
mem[1611] = 80'h0010ffabffabffabffab;
mem[1612] = 80'h0010ffabffabffabffab;
mem[1613] = 80'h0010ffabffabffabffab;
mem[1614] = 80'h0010ffabffabffabffab;
mem[1615] = 80'h0010ffabffabffabffab;
mem[1616] = 80'h0010ffabffabffabffab;
mem[1617] = 80'h0010ffabffabffabffab;
mem[1618] = 80'h0010ffabffabffabffab;
mem[1619] = 80'h0010ffabffabffabffab;
mem[1620] = 80'h0010ffabffabffabffab;
mem[1621] = 80'h0010ffabffabffabffab;
mem[1622] = 80'h0010ffabffabffabffab;
mem[1623] = 80'h0010ffabffabffabffab;
mem[1624] = 80'h0010ffabffabffabffab;
mem[1625] = 80'h0010ffabffabffabffab;
mem[1626] = 80'h0010ffabffabffabffab;
mem[1627] = 80'h0010ffabffabffabffab;
mem[1628] = 80'h0010ffabffabffabffab;
mem[1629] = 80'h0010ffabffabffabffab;
mem[1630] = 80'h0010ffabffabffabffab;
mem[1631] = 80'h0010ffabffabffabffab;
mem[1632] = 80'h0010ffabffabffabffab;
mem[1633] = 80'h0010ffabffabffabffab;
mem[1634] = 80'h0010ffabffabffabffab;
mem[1635] = 80'h0010ffabffabffabffab;
mem[1636] = 80'h0010551ac7096dc4b705;
mem[1637] = 80'h00104a192b0cdd12dd2d;
mem[1638] = 80'h011040294f822ed923b9;
mem[1639] = 80'h00000000000000000000;
mem[1640] = 80'h00000000000000000000;
mem[1641] = 80'h00000000000000000000;
mem[1642] = 80'h00000000000000000000;
mem[1643] = 80'h00000000000000000000;
mem[1644] = 80'h00000000000000000000;
mem[1645] = 80'h00000000000000000000;
mem[1646] = 80'h00000000000000000000;
mem[1647] = 80'h00000000000000000000;
mem[1648] = 80'h00000000000000000000;
mem[1649] = 80'h00000000000000000000;
mem[1650] = 80'h00000000000000000000;
mem[1651] = 80'h00000000000000000000;
mem[1652] = 80'h10100000010000010010;
mem[1653] = 80'h00109400000208004500;
mem[1654] = 80'h0010058589ab0000fffd;
mem[1655] = 80'h0010aa77c0550102c000;
mem[1656] = 80'h00100001ffabffabffab;
mem[1657] = 80'h0010ffabffabffabffab;
mem[1658] = 80'h0010ffabffabffabffab;
mem[1659] = 80'h0010ffabffabffabffab;
mem[1660] = 80'h0010ffabffabffabffab;
mem[1661] = 80'h0010ffabffabffabffab;
mem[1662] = 80'h0010ffabffabffabffab;
mem[1663] = 80'h0010ffabffabffabffab;
mem[1664] = 80'h0010ffabffabffabffab;
mem[1665] = 80'h0010ffabffabffabffab;
mem[1666] = 80'h0010ffabffabffabffab;
mem[1667] = 80'h0010ffabffabffabffab;
mem[1668] = 80'h0010ffabffabffabffab;
mem[1669] = 80'h0010ffabffabffabffab;
mem[1670] = 80'h0010ffabffabffabffab;
mem[1671] = 80'h0010ffabffabffabffab;
mem[1672] = 80'h0010ffabffabffabffab;
mem[1673] = 80'h0010ffabffabffabffab;
mem[1674] = 80'h0010ffabffabffabffab;
mem[1675] = 80'h0010ffabffabffabffab;
mem[1676] = 80'h0010ffabffabffabffab;
mem[1677] = 80'h0010ffabffabffabffab;
mem[1678] = 80'h0010ffabffabffabffab;
mem[1679] = 80'h0010ffabffabffabffab;
mem[1680] = 80'h0010ffabffabffabffab;
mem[1681] = 80'h0010ffabffabffabffab;
mem[1682] = 80'h0010ffabffabffabffab;
mem[1683] = 80'h0010ffabffabffabffab;
mem[1684] = 80'h0010ffabffabffabffab;
mem[1685] = 80'h0010ffabffabffabffab;
mem[1686] = 80'h0010ffabffabffabffab;
mem[1687] = 80'h0010ffabffabffabffab;
mem[1688] = 80'h0010ffabffabffabffab;
mem[1689] = 80'h0010ffabffabffabffab;
mem[1690] = 80'h0010ffabffabffabffab;
mem[1691] = 80'h0010ffabffabffabffab;
mem[1692] = 80'h0010ffabffabffabffab;
mem[1693] = 80'h0010ffabffabffabffab;
mem[1694] = 80'h0010ffabffabffabffab;
mem[1695] = 80'h0010ffabffabffabffab;
mem[1696] = 80'h0010ffabffabffabffab;
mem[1697] = 80'h0010ffabffabffabffab;
mem[1698] = 80'h0010ffabffabffabffab;
mem[1699] = 80'h0010ffabffabffabffab;
mem[1700] = 80'h0010ffabffabffabffab;
mem[1701] = 80'h0010ffabffabffabffab;
mem[1702] = 80'h0010ffabffabffabffab;
mem[1703] = 80'h0010ffabffabffabffab;
mem[1704] = 80'h0010ffabffabffabffab;
mem[1705] = 80'h0010ffabffabffabffab;
mem[1706] = 80'h0010ffabffabffabffab;
mem[1707] = 80'h0010ffabffabffabffab;
mem[1708] = 80'h0010ffabffabffabffab;
mem[1709] = 80'h0010ffabffabffabffab;
mem[1710] = 80'h0010ffabffabffabffab;
mem[1711] = 80'h0010ffabffabffabffab;
mem[1712] = 80'h0010ffabffabffabffab;
mem[1713] = 80'h0010ffabffabffabffab;
mem[1714] = 80'h0010ffabffabffabffab;
mem[1715] = 80'h0010ffabffabffabffab;
mem[1716] = 80'h0010ffabffabffabffab;
mem[1717] = 80'h0010ffabffabffabffab;
mem[1718] = 80'h0010ffabffabffabffab;
mem[1719] = 80'h0010ffabffabffabffab;
mem[1720] = 80'h0010ffabffabffabffab;
mem[1721] = 80'h0010ffabffabffabffab;
mem[1722] = 80'h0010ffabffabffabffab;
mem[1723] = 80'h0010ffabffabffabffab;
mem[1724] = 80'h0010ffabffabffabffab;
mem[1725] = 80'h0010ffabffabffabffab;
mem[1726] = 80'h0010ffabffabffabffab;
mem[1727] = 80'h0010ffabffabffabffab;
mem[1728] = 80'h0010ffabffabffabffab;
mem[1729] = 80'h0010ffabffabffabffab;
mem[1730] = 80'h0010ffabffabffabffab;
mem[1731] = 80'h0010ffabffabffabffab;
mem[1732] = 80'h0010ffabffabffabffab;
mem[1733] = 80'h0010ffabffabffabffab;
mem[1734] = 80'h0010ffabffabffabffab;
mem[1735] = 80'h0010ffabffabffabffab;
mem[1736] = 80'h0010ffabffabffabffab;
mem[1737] = 80'h0010ffabffabffabffab;
mem[1738] = 80'h0010ffabffabffabffab;
mem[1739] = 80'h0010ffabffabffabffab;
mem[1740] = 80'h0010ffabffabffabffab;
mem[1741] = 80'h0010ffabffabffabffab;
mem[1742] = 80'h0010ffabffabffabffab;
mem[1743] = 80'h0010ffabffabffabffab;
mem[1744] = 80'h0010ffabffabffabffab;
mem[1745] = 80'h0010ffabffabffabffab;
mem[1746] = 80'h0010ffabffabffabffab;
mem[1747] = 80'h0010ffabffabffabffab;
mem[1748] = 80'h0010ffabffabffabffab;
mem[1749] = 80'h0010ffabffabffabffab;
mem[1750] = 80'h0010ffabffabffabffab;
mem[1751] = 80'h0010ffabffabffabffab;
mem[1752] = 80'h0010ffabffabffabffab;
mem[1753] = 80'h0010ffabffabffabffab;
mem[1754] = 80'h0010ffabffabffabffab;
mem[1755] = 80'h0010ffabffabffabffab;
mem[1756] = 80'h0010ffabffabffabffab;
mem[1757] = 80'h0010ffabffabffabffab;
mem[1758] = 80'h0010ffabffabffabffab;
mem[1759] = 80'h0010ffabffabffabffab;
mem[1760] = 80'h0010ffabffabffabffab;
mem[1761] = 80'h0010ffabffabffabffab;
mem[1762] = 80'h0010ffabffabffabffab;
mem[1763] = 80'h0010ffabffabffabffab;
mem[1764] = 80'h0010ffabffabffabffab;
mem[1765] = 80'h0010ffabffabffabffab;
mem[1766] = 80'h0010ffabffabffabffab;
mem[1767] = 80'h0010ffabffabffabffab;
mem[1768] = 80'h0010ffabffabffabffab;
mem[1769] = 80'h0010ffabffabffabffab;
mem[1770] = 80'h0010ffabffabffabffab;
mem[1771] = 80'h0010ffabffabffabffab;
mem[1772] = 80'h0010ffabffabffabffab;
mem[1773] = 80'h0010ffabffabffabffab;
mem[1774] = 80'h0010ffabffabffabffab;
mem[1775] = 80'h0010ffabffabffabffab;
mem[1776] = 80'h0010ffabffabffabffab;
mem[1777] = 80'h0010ffabffabffabffab;
mem[1778] = 80'h0010ffabffabffabffab;
mem[1779] = 80'h0010ffabffabffabffab;
mem[1780] = 80'h0010ffabffabffabffab;
mem[1781] = 80'h0010ffabffabffabffab;
mem[1782] = 80'h0010ffabffabffabffab;
mem[1783] = 80'h0010ffabffabffabffab;
mem[1784] = 80'h0010ffabffabffabffab;
mem[1785] = 80'h0010ffabffabffabffab;
mem[1786] = 80'h0010ffabffabffabffab;
mem[1787] = 80'h0010ffabffabffabffab;
mem[1788] = 80'h0010ffabffabffabffab;
mem[1789] = 80'h0010ffabffabffabffab;
mem[1790] = 80'h0010ffabffabffabffab;
mem[1791] = 80'h0010ffabffabffabffab;
mem[1792] = 80'h0010ffabffabffabffab;
mem[1793] = 80'h0010ffabffabffabffab;
mem[1794] = 80'h0010ffabffabffabffab;
mem[1795] = 80'h0010ffabffabffabffab;
mem[1796] = 80'h0010ffabffabffabffab;
mem[1797] = 80'h0010ffabffabffabffab;
mem[1798] = 80'h0010ffabffabffabffab;
mem[1799] = 80'h0010ffabffabffabffab;
mem[1800] = 80'h0010ffabffabffabffab;
mem[1801] = 80'h0010ffabffabffabffab;
mem[1802] = 80'h0010ffabffabffabffab;
mem[1803] = 80'h0010ffabffabffabffab;
mem[1804] = 80'h0010ffabffabffabffab;
mem[1805] = 80'h0010ffabffabffabffab;
mem[1806] = 80'h0010ffabffabffabffab;
mem[1807] = 80'h0010ffabffabffabffab;
mem[1808] = 80'h0010ffabffabffabffab;
mem[1809] = 80'h0010ffabffabffabffab;
mem[1810] = 80'h0010ffabffabffabffab;
mem[1811] = 80'h0010ffabffabffabffab;
mem[1812] = 80'h0010ffabffabffabffab;
mem[1813] = 80'h0010ffabffabffabffab;
mem[1814] = 80'h0010ffabffabffabffab;
mem[1815] = 80'h0010ffabffabffabffab;
mem[1816] = 80'h0010ffabffabffabffab;
mem[1817] = 80'h0010ffabffabffabffab;
mem[1818] = 80'h0010ffabffabffabffab;
mem[1819] = 80'h0010ffabffabffabffab;
mem[1820] = 80'h0010ffabffabffabffab;
mem[1821] = 80'h0010ffabffabffabffab;
mem[1822] = 80'h0010ffabffabffabffab;
mem[1823] = 80'h0010ffabffabffabffab;
mem[1824] = 80'h0010ffabffabffabffab;
mem[1825] = 80'h0010ffabffabffabffab;
mem[1826] = 80'h0010ffabffabffabffab;
mem[1827] = 80'h0010ffabffabffabff54;
mem[1828] = 80'h00106b1925b5bd75ba81;
mem[1829] = 80'h0010cbace128c0cf7c3a;
mem[1830] = 80'h011792057b841cefa200;
mem[1831] = 80'h00000000000000000000;
mem[1832] = 80'h00000000000000000000;
mem[1833] = 80'h00000000000000000000;
mem[1834] = 80'h00000000000000000000;
mem[1835] = 80'h00000000000000000000;
mem[1836] = 80'h00000000000000000000;
mem[1837] = 80'h00000000000000000000;
mem[1838] = 80'h00000000000000000000;
mem[1839] = 80'h10100000010000010010;
mem[1840] = 80'h00109400000208004500;
mem[1841] = 80'h001005af89ac0000fffd;
mem[1842] = 80'h0010aa4cc0550102c000;
mem[1843] = 80'h00100001ffabffabffab;
mem[1844] = 80'h0010ffabffabffabffab;
mem[1845] = 80'h0010ffabffabffabffab;
mem[1846] = 80'h0010ffabffabffabffab;
mem[1847] = 80'h0010ffabffabffabffab;
mem[1848] = 80'h0010ffabffabffabffab;
mem[1849] = 80'h0010ffabffabffabffab;
mem[1850] = 80'h0010ffabffabffabffab;
mem[1851] = 80'h0010ffabffabffabffab;
mem[1852] = 80'h0010ffabffabffabffab;
mem[1853] = 80'h0010ffabffabffabffab;
mem[1854] = 80'h0010ffabffabffabffab;
mem[1855] = 80'h0010ffabffabffabffab;
mem[1856] = 80'h0010ffabffabffabffab;
mem[1857] = 80'h0010ffabffabffabffab;
mem[1858] = 80'h0010ffabffabffabffab;
mem[1859] = 80'h0010ffabffabffabffab;
mem[1860] = 80'h0010ffabffabffabffab;
mem[1861] = 80'h0010ffabffabffabffab;
mem[1862] = 80'h0010ffabffabffabffab;
mem[1863] = 80'h0010ffabffabffabffab;
mem[1864] = 80'h0010ffabffabffabffab;
mem[1865] = 80'h0010ffabffabffabffab;
mem[1866] = 80'h0010ffabffabffabffab;
mem[1867] = 80'h0010ffabffabffabffab;
mem[1868] = 80'h0010ffabffabffabffab;
mem[1869] = 80'h0010ffabffabffabffab;
mem[1870] = 80'h0010ffabffabffabffab;
mem[1871] = 80'h0010ffabffabffabffab;
mem[1872] = 80'h0010ffabffabffabffab;
mem[1873] = 80'h0010ffabffabffabffab;
mem[1874] = 80'h0010ffabffabffabffab;
mem[1875] = 80'h0010ffabffabffabffab;
mem[1876] = 80'h0010ffabffabffabffab;
mem[1877] = 80'h0010ffabffabffabffab;
mem[1878] = 80'h0010ffabffabffabffab;
mem[1879] = 80'h0010ffabffabffabffab;
mem[1880] = 80'h0010ffabffabffabffab;
mem[1881] = 80'h0010ffabffabffabffab;
mem[1882] = 80'h0010ffabffabffabffab;
mem[1883] = 80'h0010ffabffabffabffab;
mem[1884] = 80'h0010ffabffabffabffab;
mem[1885] = 80'h0010ffabffabffabffab;
mem[1886] = 80'h0010ffabffabffabffab;
mem[1887] = 80'h0010ffabffabffabffab;
mem[1888] = 80'h0010ffabffabffabffab;
mem[1889] = 80'h0010ffabffabffabffab;
mem[1890] = 80'h0010ffabffabffabffab;
mem[1891] = 80'h0010ffabffabffabffab;
mem[1892] = 80'h0010ffabffabffabffab;
mem[1893] = 80'h0010ffabffabffabffab;
mem[1894] = 80'h0010ffabffabffabffab;
mem[1895] = 80'h0010ffabffabffabffab;
mem[1896] = 80'h0010ffabffabffabffab;
mem[1897] = 80'h0010ffabffabffabffab;
mem[1898] = 80'h0010ffabffabffabffab;
mem[1899] = 80'h0010ffabffabffabffab;
mem[1900] = 80'h0010ffabffabffabffab;
mem[1901] = 80'h0010ffabffabffabffab;
mem[1902] = 80'h0010ffabffabffabffab;
mem[1903] = 80'h0010ffabffabffabffab;
mem[1904] = 80'h0010ffabffabffabffab;
mem[1905] = 80'h0010ffabffabffabffab;
mem[1906] = 80'h0010ffabffabffabffab;
mem[1907] = 80'h0010ffabffabffabffab;
mem[1908] = 80'h0010ffabffabffabffab;
mem[1909] = 80'h0010ffabffabffabffab;
mem[1910] = 80'h0010ffabffabffabffab;
mem[1911] = 80'h0010ffabffabffabffab;
mem[1912] = 80'h0010ffabffabffabffab;
mem[1913] = 80'h0010ffabffabffabffab;
mem[1914] = 80'h0010ffabffabffabffab;
mem[1915] = 80'h0010ffabffabffabffab;
mem[1916] = 80'h0010ffabffabffabffab;
mem[1917] = 80'h0010ffabffabffabffab;
mem[1918] = 80'h0010ffabffabffabffab;
mem[1919] = 80'h0010ffabffabffabffab;
mem[1920] = 80'h0010ffabffabffabffab;
mem[1921] = 80'h0010ffabffabffabffab;
mem[1922] = 80'h0010ffabffabffabffab;
mem[1923] = 80'h0010ffabffabffabffab;
mem[1924] = 80'h0010ffabffabffabffab;
mem[1925] = 80'h0010ffabffabffabffab;
mem[1926] = 80'h0010ffabffabffabffab;
mem[1927] = 80'h0010ffabffabffabffab;
mem[1928] = 80'h0010ffabffabffabffab;
mem[1929] = 80'h0010ffabffabffabffab;
mem[1930] = 80'h0010ffabffabffabffab;
mem[1931] = 80'h0010ffabffabffabffab;
mem[1932] = 80'h0010ffabffabffabffab;
mem[1933] = 80'h0010ffabffabffabffab;
mem[1934] = 80'h0010ffabffabffabffab;
mem[1935] = 80'h0010ffabffabffabffab;
mem[1936] = 80'h0010ffabffabffabffab;
mem[1937] = 80'h0010ffabffabffabffab;
mem[1938] = 80'h0010ffabffabffabffab;
mem[1939] = 80'h0010ffabffabffabffab;
mem[1940] = 80'h0010ffabffabffabffab;
mem[1941] = 80'h0010ffabffabffabffab;
mem[1942] = 80'h0010ffabffabffabffab;
mem[1943] = 80'h0010ffabffabffabffab;
mem[1944] = 80'h0010ffabffabffabffab;
mem[1945] = 80'h0010ffabffabffabffab;
mem[1946] = 80'h0010ffabffabffabffab;
mem[1947] = 80'h0010ffabffabffabffab;
mem[1948] = 80'h0010ffabffabffabffab;
mem[1949] = 80'h0010ffabffabffabffab;
mem[1950] = 80'h0010ffabffabffabffab;
mem[1951] = 80'h0010ffabffabffabffab;
mem[1952] = 80'h0010ffabffabffabffab;
mem[1953] = 80'h0010ffabffabffabffab;
mem[1954] = 80'h0010ffabffabffabffab;
mem[1955] = 80'h0010ffabffabffabffab;
mem[1956] = 80'h0010ffabffabffabffab;
mem[1957] = 80'h0010ffabffabffabffab;
mem[1958] = 80'h0010ffabffabffabffab;
mem[1959] = 80'h0010ffabffabffabffab;
mem[1960] = 80'h0010ffabffabffabffab;
mem[1961] = 80'h0010ffabffabffabffab;
mem[1962] = 80'h0010ffabffabffabffab;
mem[1963] = 80'h0010ffabffabffabffab;
mem[1964] = 80'h0010ffabffabffabffab;
mem[1965] = 80'h0010ffabffabffabffab;
mem[1966] = 80'h0010ffabffabffabffab;
mem[1967] = 80'h0010ffabffabffabffab;
mem[1968] = 80'h0010ffabffabffabffab;
mem[1969] = 80'h0010ffabffabffabffab;
mem[1970] = 80'h0010ffabffabffabffab;
mem[1971] = 80'h0010ffabffabffabffab;
mem[1972] = 80'h0010ffabffabffabffab;
mem[1973] = 80'h0010ffabffabffabffab;
mem[1974] = 80'h0010ffabffabffabffab;
mem[1975] = 80'h0010ffabffabffabffab;
mem[1976] = 80'h0010ffabffabffabffab;
mem[1977] = 80'h0010ffabffabffabffab;
mem[1978] = 80'h0010ffabffabffabffab;
mem[1979] = 80'h0010ffabffabffabffab;
mem[1980] = 80'h0010ffabffabffabffab;
mem[1981] = 80'h0010ffabffabffabffab;
mem[1982] = 80'h0010ffabffabffabffab;
mem[1983] = 80'h0010ffabffabffabffab;
mem[1984] = 80'h0010ffabffabffabffab;
mem[1985] = 80'h0010ffabffabffabffab;
mem[1986] = 80'h0010ffabffabffabffab;
mem[1987] = 80'h0010ffabffabffabffab;
mem[1988] = 80'h0010ffabffabffabffab;
mem[1989] = 80'h0010ffabffabffabffab;
mem[1990] = 80'h0010ffabffabffabffab;
mem[1991] = 80'h0010ffabffabffabffab;
mem[1992] = 80'h0010ffabffabffabffab;
mem[1993] = 80'h0010ffabffabffabffab;
mem[1994] = 80'h0010ffabffabffabffab;
mem[1995] = 80'h0010ffabffabffabffab;
mem[1996] = 80'h0010ffabffabffabffab;
mem[1997] = 80'h0010ffabffabffabffab;
mem[1998] = 80'h0010ffabffabffabffab;
mem[1999] = 80'h0010ffabffabffabffab;
mem[2000] = 80'h0010ffabffabffabffab;
mem[2001] = 80'h0010ffabffabffabffab;
mem[2002] = 80'h0010ffabffabffabffab;
mem[2003] = 80'h0010ffabffabffabffab;
mem[2004] = 80'h0010ffabffabffabffab;
mem[2005] = 80'h0010ffabffabffabffab;
mem[2006] = 80'h0010ffabffabffabffab;
mem[2007] = 80'h0010ffabffabffabffab;
mem[2008] = 80'h0010ffabffabffabffab;
mem[2009] = 80'h0010ffabffabffabffab;
mem[2010] = 80'h0010ffabffabffabffab;
mem[2011] = 80'h0010ffabffabffabffab;
mem[2012] = 80'h0010ffabffabffabffab;
mem[2013] = 80'h0010ffabffabffabffab;
mem[2014] = 80'h0010ffabffabffabffab;
mem[2015] = 80'h0010ffabffabffabffab;
mem[2016] = 80'h0010ffabffabffabffab;
mem[2017] = 80'h0010ffabffabffabffab;
mem[2018] = 80'h0010ffabffabffabffab;
mem[2019] = 80'h0010ffabffabffabffab;
mem[2020] = 80'h0010ff534fddcf64a9fa;
mem[2021] = 80'h00103a3924bd8d142060;
mem[2022] = 80'h00109945bdbed3be9ef8;
mem[2023] = 80'h01119300000000000000;
mem[2024] = 80'h10100000010000010010;
mem[2025] = 80'h00109400000208004500;
mem[2026] = 80'h001002ee89ad0000fffd;
mem[2027] = 80'h0010ad0cc0550102c000;
mem[2028] = 80'h00100001ffabffabffab;
mem[2029] = 80'h0010ffabffabffabffab;
mem[2030] = 80'h0010ffabffabffabffab;
mem[2031] = 80'h0010ffabffabffabffab;
mem[2032] = 80'h0010ffabffabffabffab;
mem[2033] = 80'h0010ffabffabffabffab;
mem[2034] = 80'h0010ffabffabffabffab;
mem[2035] = 80'h0010ffabffabffabffab;
mem[2036] = 80'h0010ffabffabffabffab;
mem[2037] = 80'h0010ffabffabffabffab;
mem[2038] = 80'h0010ffabffabffabffab;
mem[2039] = 80'h0010ffabffabffabffab;
mem[2040] = 80'h0010ffabffabffabffab;
mem[2041] = 80'h0010ffabffabffabffab;
mem[2042] = 80'h0010ffabffabffabffab;
mem[2043] = 80'h0010ffabffabffabffab;
mem[2044] = 80'h0010ffabffabffabffab;
mem[2045] = 80'h0010ffabffabffabffab;
mem[2046] = 80'h0010ffabffabffabffab;
mem[2047] = 80'h0010ffabffabffabffab;
mem[2048] = 80'h0010ffabffabffabffab;
mem[2049] = 80'h0010ffabffabffabffab;
mem[2050] = 80'h0010ffabffabffabffab;
mem[2051] = 80'h0010ffabffabffabffab;
mem[2052] = 80'h0010ffabffabffabffab;
mem[2053] = 80'h0010ffabffabffabffab;
mem[2054] = 80'h0010ffabffabffabffab;
mem[2055] = 80'h0010ffabffabffabffab;
mem[2056] = 80'h0010ffabffabffabffab;
mem[2057] = 80'h0010ffabffabffabffab;
mem[2058] = 80'h0010ffabffabffabffab;
mem[2059] = 80'h0010ffabffabffabffab;
mem[2060] = 80'h0010ffabffabffabffab;
mem[2061] = 80'h0010ffabffabffabffab;
mem[2062] = 80'h0010ffabffabffabffab;
mem[2063] = 80'h0010ffabffabffabffab;
mem[2064] = 80'h0010ffabffabffabffab;
mem[2065] = 80'h0010ffabffabffabffab;
mem[2066] = 80'h0010ffabffabffabffab;
mem[2067] = 80'h0010ffabffabffabffab;
mem[2068] = 80'h0010ffabffabffabffab;
mem[2069] = 80'h0010ffabffabffabffab;
mem[2070] = 80'h0010ffabffabffabffab;
mem[2071] = 80'h0010ffabffabffabffab;
mem[2072] = 80'h0010ffabffabffabffab;
mem[2073] = 80'h0010ffabffabffabffab;
mem[2074] = 80'h0010ffabffabffabffab;
mem[2075] = 80'h0010ffabffabffabffab;
mem[2076] = 80'h0010ffabffabffabffab;
mem[2077] = 80'h0010ffabffabffabffab;
mem[2078] = 80'h0010ffabffabffabffab;
mem[2079] = 80'h0010ffabffabffabffab;
mem[2080] = 80'h0010ffabffabffabffab;
mem[2081] = 80'h0010ffabffabffabffab;
mem[2082] = 80'h0010ffabffabffabffab;
mem[2083] = 80'h0010ffabffabffabffab;
mem[2084] = 80'h0010ffabffabffabffab;
mem[2085] = 80'h0010ffabffabffabffab;
mem[2086] = 80'h0010ffabffabffabffab;
mem[2087] = 80'h0010ffabffabffabffab;
mem[2088] = 80'h0010ffabffabffabffab;
mem[2089] = 80'h0010ffabffabffabffab;
mem[2090] = 80'h0010ffabffabffabffab;
mem[2091] = 80'h0010ffabffabffabffab;
mem[2092] = 80'h0010ffabffabffabffab;
mem[2093] = 80'h0010ffabffabffabffab;
mem[2094] = 80'h0010ffabffabffabffab;
mem[2095] = 80'h0010ffabffabffabffab;
mem[2096] = 80'h0010ffabffabffabffab;
mem[2097] = 80'h0010ffabffabffabffab;
mem[2098] = 80'h0010ffabffabffabffab;
mem[2099] = 80'h0010ffabffabffabffab;
mem[2100] = 80'h0010ffabffabffabffab;
mem[2101] = 80'h0010ffabffabffabffab;
mem[2102] = 80'h0010ffabffabffabffab;
mem[2103] = 80'h0010ffabffabffabffab;
mem[2104] = 80'h0010ffabffabffabffab;
mem[2105] = 80'h0010ffabffabffabffab;
mem[2106] = 80'h0010ffabffabffabffab;
mem[2107] = 80'h0010ffabffabffabffab;
mem[2108] = 80'h0010ffabffabffabffab;
mem[2109] = 80'h0010ffabffabffabffab;
mem[2110] = 80'h0010ffabffabffabffab;
mem[2111] = 80'h0010ffabffabffabffab;
mem[2112] = 80'h0010ffabffabffabffab;
mem[2113] = 80'h0010ffabffabffabffab;
mem[2114] = 80'h0010ffabffabffabffab;
mem[2115] = 80'h0010ffabffabffabffab;
mem[2116] = 80'h0010ffabffabffabffab;
mem[2117] = 80'h0010523e03e3bcd03885;
mem[2118] = 80'h0010f2f63a60e1f627c8;
mem[2119] = 80'h0110128c6ae6e797baa8;
mem[2120] = 80'h10100000010000010010;
mem[2121] = 80'h00109400000208004500;
mem[2122] = 80'h0010018e89ae0000fffd;
mem[2123] = 80'h0010ae6bc0550102c000;
mem[2124] = 80'h00100001ffabffabffab;
mem[2125] = 80'h0010ffabffabffabffab;
mem[2126] = 80'h0010ffabffabffabffab;
mem[2127] = 80'h0010ffabffabffabffab;
mem[2128] = 80'h0010ffabffabffabffab;
mem[2129] = 80'h0010ffabffabffabffab;
mem[2130] = 80'h0010ffabffabffabffab;
mem[2131] = 80'h0010ffabffabffabffab;
mem[2132] = 80'h0010ffabffabffabffab;
mem[2133] = 80'h0010ffabffabffabffab;
mem[2134] = 80'h0010ffabffabffabffab;
mem[2135] = 80'h0010ffabffabffabffab;
mem[2136] = 80'h0010ffabffabffabffab;
mem[2137] = 80'h0010ffabffabffabffab;
mem[2138] = 80'h0010ffabffabffabffab;
mem[2139] = 80'h0010ffabffabffabffab;
mem[2140] = 80'h0010ffabffabffabffab;
mem[2141] = 80'h0010ffabffabffabffab;
mem[2142] = 80'h0010ffabffabffabffab;
mem[2143] = 80'h0010ffabffabffabffab;
mem[2144] = 80'h0010ffabffabffabffab;
mem[2145] = 80'h0010ffabffabffabffab;
mem[2146] = 80'h0010ffabffabffabffab;
mem[2147] = 80'h0010ffabffabffabffab;
mem[2148] = 80'h0010ffabffabffabffab;
mem[2149] = 80'h0010ffabffabffabffab;
mem[2150] = 80'h0010ffabffabffabffab;
mem[2151] = 80'h0010ffabffabffabffab;
mem[2152] = 80'h0010ffabffabffabffab;
mem[2153] = 80'h0010ffabffabffabffab;
mem[2154] = 80'h0010ffabffabffabffab;
mem[2155] = 80'h0010ffabffabffabffab;
mem[2156] = 80'h0010ffabffabffabffab;
mem[2157] = 80'h0010ffabffabffabffab;
mem[2158] = 80'h0010ffabffabffabffab;
mem[2159] = 80'h0010ffabffabffabffab;
mem[2160] = 80'h0010ffabffabffabffab;
mem[2161] = 80'h0010ffabffabffabffab;
mem[2162] = 80'h0010ffabffabffabffab;
mem[2163] = 80'h0010ffabffabffabffab;
mem[2164] = 80'h0010ffabffabffabffab;
mem[2165] = 80'h0010ffabffabffabffab;
mem[2166] = 80'h0010ffabffabffabffab;
mem[2167] = 80'h0010ffabffabffabffab;
mem[2168] = 80'h0010ffabffabffabffab;
mem[2169] = 80'h001051ac6196d45a7f45;
mem[2170] = 80'h0010ae81b256ff858e3a;
mem[2171] = 80'h01106e459c3ed7ddd217;
mem[2172] = 80'h10100000010000010010;
mem[2173] = 80'h00109400000208004500;
mem[2174] = 80'h001003b789af0000fffd;
mem[2175] = 80'h0010ac41c0550102c000;
mem[2176] = 80'h00100001ffabffabffab;
mem[2177] = 80'h0010ffabffabffabffab;
mem[2178] = 80'h0010ffabffabffabffab;
mem[2179] = 80'h0010ffabffabffabffab;
mem[2180] = 80'h0010ffabffabffabffab;
mem[2181] = 80'h0010ffabffabffabffab;
mem[2182] = 80'h0010ffabffabffabffab;
mem[2183] = 80'h0010ffabffabffabffab;
mem[2184] = 80'h0010ffabffabffabffab;
mem[2185] = 80'h0010ffabffabffabffab;
mem[2186] = 80'h0010ffabffabffabffab;
mem[2187] = 80'h0010ffabffabffabffab;
mem[2188] = 80'h0010ffabffabffabffab;
mem[2189] = 80'h0010ffabffabffabffab;
mem[2190] = 80'h0010ffabffabffabffab;
mem[2191] = 80'h0010ffabffabffabffab;
mem[2192] = 80'h0010ffabffabffabffab;
mem[2193] = 80'h0010ffabffabffabffab;
mem[2194] = 80'h0010ffabffabffabffab;
mem[2195] = 80'h0010ffabffabffabffab;
mem[2196] = 80'h0010ffabffabffabffab;
mem[2197] = 80'h0010ffabffabffabffab;
mem[2198] = 80'h0010ffabffabffabffab;
mem[2199] = 80'h0010ffabffabffabffab;
mem[2200] = 80'h0010ffabffabffabffab;
mem[2201] = 80'h0010ffabffabffabffab;
mem[2202] = 80'h0010ffabffabffabffab;
mem[2203] = 80'h0010ffabffabffabffab;
mem[2204] = 80'h0010ffabffabffabffab;
mem[2205] = 80'h0010ffabffabffabffab;
mem[2206] = 80'h0010ffabffabffabffab;
mem[2207] = 80'h0010ffabffabffabffab;
mem[2208] = 80'h0010ffabffabffabffab;
mem[2209] = 80'h0010ffabffabffabffab;
mem[2210] = 80'h0010ffabffabffabffab;
mem[2211] = 80'h0010ffabffabffabffab;
mem[2212] = 80'h0010ffabffabffabffab;
mem[2213] = 80'h0010ffabffabffabffab;
mem[2214] = 80'h0010ffabffabffabffab;
mem[2215] = 80'h0010ffabffabffabffab;
mem[2216] = 80'h0010ffabffabffabffab;
mem[2217] = 80'h0010ffabffabffabffab;
mem[2218] = 80'h0010ffabffabffabffab;
mem[2219] = 80'h0010ffabffabffabffab;
mem[2220] = 80'h0010ffabffabffabffab;
mem[2221] = 80'h0010ffabffabffabffab;
mem[2222] = 80'h0010ffabffabffabffab;
mem[2223] = 80'h0010ffabffabffabffab;
mem[2224] = 80'h0010ffabffabffabffab;
mem[2225] = 80'h0010ffabffabffabffab;
mem[2226] = 80'h0010ffabffabffabffab;
mem[2227] = 80'h0010ffabffabffabffab;
mem[2228] = 80'h0010ffabffabffabffab;
mem[2229] = 80'h0010ffabffabffabffab;
mem[2230] = 80'h0010ffabffabffabffab;
mem[2231] = 80'h0010ffabffabffabffab;
mem[2232] = 80'h0010ffabffabffabffab;
mem[2233] = 80'h0010ffabffabffabffab;
mem[2234] = 80'h0010ffabffabffabffab;
mem[2235] = 80'h0010ffabffabffabffab;
mem[2236] = 80'h0010ffabffabffabffab;
mem[2237] = 80'h0010ffabffabffabffab;
mem[2238] = 80'h0010ffabffabffabffab;
mem[2239] = 80'h0010ffabffabffabffab;
mem[2240] = 80'h0010ffabffabffabffab;
mem[2241] = 80'h0010ffabffabffabffab;
mem[2242] = 80'h0010ffabffabffabffab;
mem[2243] = 80'h0010ffabffabffabffab;
mem[2244] = 80'h0010ffabffabffabffab;
mem[2245] = 80'h0010ffabffabffabffab;
mem[2246] = 80'h0010ffabffabffabffab;
mem[2247] = 80'h0010ffabffabffabffab;
mem[2248] = 80'h0010ffabffabffabffab;
mem[2249] = 80'h0010ffabffabffabffab;
mem[2250] = 80'h0010ffabffabffabffab;
mem[2251] = 80'h0010ffabffabffabffab;
mem[2252] = 80'h0010ffabffabffabffab;
mem[2253] = 80'h0010ffabffabffabffab;
mem[2254] = 80'h0010ffabffabffabffab;
mem[2255] = 80'h0010ffabffabffabffab;
mem[2256] = 80'h0010ffabffabffabffab;
mem[2257] = 80'h0010ffabffabffabffab;
mem[2258] = 80'h0010ffabffabffabffab;
mem[2259] = 80'h0010ffabffabffabffab;
mem[2260] = 80'h0010ffabffabffabffab;
mem[2261] = 80'h0010ffabffabffabffab;
mem[2262] = 80'h0010ffabffabffabffab;
mem[2263] = 80'h0010ffabffabffabffab;
mem[2264] = 80'h0010ffabffabffabffab;
mem[2265] = 80'h0010ffabffabffabffab;
mem[2266] = 80'h0010ffabffabffabffab;
mem[2267] = 80'h0010ffabffabffabffab;
mem[2268] = 80'h0010ffabffabffabffab;
mem[2269] = 80'h0010ffabffabffabffab;
mem[2270] = 80'h0010ffabffabffabffab;
mem[2271] = 80'h0010ffabffabffabffab;
mem[2272] = 80'h0010ffabffabffabffab;
mem[2273] = 80'h0010ffabffabffabffab;
mem[2274] = 80'h0010ffabffabffabffab;
mem[2275] = 80'h0010ffabffabffabffab;
mem[2276] = 80'h0010ffabffabffabffab;
mem[2277] = 80'h0010ffabffabffabffab;
mem[2278] = 80'h0010ffabffabffabffab;
mem[2279] = 80'h0010ffabffabffabffab;
mem[2280] = 80'h0010ffabffabffabffab;
mem[2281] = 80'h0010ffabffabffabffab;
mem[2282] = 80'h0010ffabffabffabffab;
mem[2283] = 80'h0010ffabffabffabffab;
mem[2284] = 80'h0010ffabffabffabffab;
mem[2285] = 80'h0010ffabffabffabffab;
mem[2286] = 80'h0010ffabffabffabffab;
mem[2287] = 80'h0010ffabffabffabffab;
mem[2288] = 80'h0010ffabffabffabffab;
mem[2289] = 80'h0010ffabffabffabffab;
mem[2290] = 80'h0010ff50ddbfba0c23bd;
mem[2291] = 80'h0010fa655335bb0a5476;
mem[2292] = 80'h00106bb2d756a452a992;
mem[2293] = 80'h0111be00000000000000;
mem[2294] = 80'h10100000010000010010;
mem[2295] = 80'h00109400000208004500;
mem[2296] = 80'h001004cb89b00000fffd;
mem[2297] = 80'h0010ab2cc0550102c000;
mem[2298] = 80'h00100001ffabffabffab;
mem[2299] = 80'h0010ffabffabffabffab;
mem[2300] = 80'h0010ffabffabffabffab;
mem[2301] = 80'h0010ffabffabffabffab;
mem[2302] = 80'h0010ffabffabffabffab;
mem[2303] = 80'h0010ffabffabffabffab;
mem[2304] = 80'h0010ffabffabffabffab;
mem[2305] = 80'h0010ffabffabffabffab;
mem[2306] = 80'h0010ffabffabffabffab;
mem[2307] = 80'h0010ffabffabffabffab;
mem[2308] = 80'h0010ffabffabffabffab;
mem[2309] = 80'h0010ffabffabffabffab;
mem[2310] = 80'h0010ffabffabffabffab;
mem[2311] = 80'h0010ffabffabffabffab;
mem[2312] = 80'h0010ffabffabffabffab;
mem[2313] = 80'h0010ffabffabffabffab;
mem[2314] = 80'h0010ffabffabffabffab;
mem[2315] = 80'h0010ffabffabffabffab;
mem[2316] = 80'h0010ffabffabffabffab;
mem[2317] = 80'h0010ffabffabffabffab;
mem[2318] = 80'h0010ffabffabffabffab;
mem[2319] = 80'h0010ffabffabffabffab;
mem[2320] = 80'h0010ffabffabffabffab;
mem[2321] = 80'h0010ffabffabffabffab;
mem[2322] = 80'h0010ffabffabffabffab;
mem[2323] = 80'h0010ffabffabffabffab;
mem[2324] = 80'h0010ffabffabffabffab;
mem[2325] = 80'h0010ffabffabffabffab;
mem[2326] = 80'h0010ffabffabffabffab;
mem[2327] = 80'h0010ffabffabffabffab;
mem[2328] = 80'h0010ffabffabffabffab;
mem[2329] = 80'h0010ffabffabffabffab;
mem[2330] = 80'h0010ffabffabffabffab;
mem[2331] = 80'h0010ffabffabffabffab;
mem[2332] = 80'h0010ffabffabffabffab;
mem[2333] = 80'h0010ffabffabffabffab;
mem[2334] = 80'h0010ffabffabffabffab;
mem[2335] = 80'h0010ffabffabffabffab;
mem[2336] = 80'h0010ffabffabffabffab;
mem[2337] = 80'h0010ffabffabffabffab;
mem[2338] = 80'h0010ffabffabffabffab;
mem[2339] = 80'h0010ffabffabffabffab;
mem[2340] = 80'h0010ffabffabffabffab;
mem[2341] = 80'h0010ffabffabffabffab;
mem[2342] = 80'h0010ffabffabffabffab;
mem[2343] = 80'h0010ffabffabffabffab;
mem[2344] = 80'h0010ffabffabffabffab;
mem[2345] = 80'h0010ffabffabffabffab;
mem[2346] = 80'h0010ffabffabffabffab;
mem[2347] = 80'h0010ffabffabffabffab;
mem[2348] = 80'h0010ffabffabffabffab;
mem[2349] = 80'h0010ffabffabffabffab;
mem[2350] = 80'h0010ffabffabffabffab;
mem[2351] = 80'h0010ffabffabffabffab;
mem[2352] = 80'h0010ffabffabffabffab;
mem[2353] = 80'h0010ffabffabffabffab;
mem[2354] = 80'h0010ffabffabffabffab;
mem[2355] = 80'h0010ffabffabffabffab;
mem[2356] = 80'h0010ffabffabffabffab;
mem[2357] = 80'h0010ffabffabffabffab;
mem[2358] = 80'h0010ffabffabffabffab;
mem[2359] = 80'h0010ffabffabffabffab;
mem[2360] = 80'h0010ffabffabffabffab;
mem[2361] = 80'h0010ffabffabffabffab;
mem[2362] = 80'h0010ffabffabffabffab;
mem[2363] = 80'h0010ffabffabffabffab;
mem[2364] = 80'h0010ffabffabffabffab;
mem[2365] = 80'h0010ffabffabffabffab;
mem[2366] = 80'h0010ffabffabffabffab;
mem[2367] = 80'h0010ffabffabffabffab;
mem[2368] = 80'h0010ffabffabffabffab;
mem[2369] = 80'h0010ffabffabffabffab;
mem[2370] = 80'h0010ffabffabffabffab;
mem[2371] = 80'h0010ffabffabffabffab;
mem[2372] = 80'h0010ffabffabffabffab;
mem[2373] = 80'h0010ffabffabffabffab;
mem[2374] = 80'h0010ffabffabffabffab;
mem[2375] = 80'h0010ffabffabffabffab;
mem[2376] = 80'h0010ffabffabffabffab;
mem[2377] = 80'h0010ffabffabffabffab;
mem[2378] = 80'h0010ffabffabffabffab;
mem[2379] = 80'h0010ffabffabffabffab;
mem[2380] = 80'h0010ffabffabffabffab;
mem[2381] = 80'h0010ffabffabffabffab;
mem[2382] = 80'h0010ffabffabffabffab;
mem[2383] = 80'h0010ffabffabffabffab;
mem[2384] = 80'h0010ffabffabffabffab;
mem[2385] = 80'h0010ffabffabffabffab;
mem[2386] = 80'h0010ffabffabffabffab;
mem[2387] = 80'h0010ffabffabffabffab;
mem[2388] = 80'h0010ffabffabffabffab;
mem[2389] = 80'h0010ffabffabffabffab;
mem[2390] = 80'h0010ffabffabffabffab;
mem[2391] = 80'h0010ffabffabffabffab;
mem[2392] = 80'h0010ffabffabffabffab;
mem[2393] = 80'h0010ffabffabffabffab;
mem[2394] = 80'h0010ffabffabffabffab;
mem[2395] = 80'h0010ffabffabffabffab;
mem[2396] = 80'h0010ffabffabffabffab;
mem[2397] = 80'h0010ffabffabffabffab;
mem[2398] = 80'h0010ffabffabffabffab;
mem[2399] = 80'h0010ffabffabffabffab;
mem[2400] = 80'h0010ffabffabffabffab;
mem[2401] = 80'h0010ffabffabffabffab;
mem[2402] = 80'h0010ffabffabffabffab;
mem[2403] = 80'h0010ffabffabffabffab;
mem[2404] = 80'h0010ffabffabffabffab;
mem[2405] = 80'h0010ffabffabffabffab;
mem[2406] = 80'h0010ffabffabffabffab;
mem[2407] = 80'h0010ffabffabffabffab;
mem[2408] = 80'h0010ffabffabffabffab;
mem[2409] = 80'h0010ffabffabffabffab;
mem[2410] = 80'h0010ffabffabffabffab;
mem[2411] = 80'h0010ffabffabffabffab;
mem[2412] = 80'h0010ffabffabffabffab;
mem[2413] = 80'h0010ffabffabffabffab;
mem[2414] = 80'h0010ffabffabffabffab;
mem[2415] = 80'h0010ffabffabffabffab;
mem[2416] = 80'h0010ffabffabffabffab;
mem[2417] = 80'h0010ffabffabffabffab;
mem[2418] = 80'h0010ffabffabffabffab;
mem[2419] = 80'h0010ffabffabffabffab;
mem[2420] = 80'h0010ffabffabffabffab;
mem[2421] = 80'h0010ffabffabffabffab;
mem[2422] = 80'h0010ffabffabffabffab;
mem[2423] = 80'h0010ffabffabffabffab;
mem[2424] = 80'h0010ffabffabffabffab;
mem[2425] = 80'h0010ffabffabffabffab;
mem[2426] = 80'h0010ffabffabffabffab;
mem[2427] = 80'h0010ffabffabffabffab;
mem[2428] = 80'h0010ffabffabffabffab;
mem[2429] = 80'h0010ffabffabffabffab;
mem[2430] = 80'h0010ffabffabffabffab;
mem[2431] = 80'h0010ffabffabffabffab;
mem[2432] = 80'h0010ffabffabffabffab;
mem[2433] = 80'h0010ffabffabffabffab;
mem[2434] = 80'h0010ffabffabffabffab;
mem[2435] = 80'h0010ffabffabffabffab;
mem[2436] = 80'h0010ffabffabffabffab;
mem[2437] = 80'h0010ffabffabffabffab;
mem[2438] = 80'h0010ffabffabffabffab;
mem[2439] = 80'h0010ffabffabffabffab;
mem[2440] = 80'h0010ffabffabffabffab;
mem[2441] = 80'h0010ffabffabffabffab;
mem[2442] = 80'h0010ffabffabffabffab;
mem[2443] = 80'h0010ffabffabffabffab;
mem[2444] = 80'h0010ffabffabffabffab;
mem[2445] = 80'h0010ffabffabffabffab;
mem[2446] = 80'h0010ffabffabff4fdcce;
mem[2447] = 80'h00106420fbc438da98f8;
mem[2448] = 80'h00103de7be650e5e877e;
mem[2449] = 80'h01155f0491c29a000000;
mem[2450] = 80'h10100000010000010010;
mem[2451] = 80'h00109400000208004500;
mem[2452] = 80'h0010027b89b10000fffd;
mem[2453] = 80'h0010ad7bc0550102c000;
mem[2454] = 80'h00100001ffabffabffab;
mem[2455] = 80'h0010ffabffabffabffab;
mem[2456] = 80'h0010ffabffabffabffab;
mem[2457] = 80'h0010ffabffabffabffab;
mem[2458] = 80'h0010ffabffabffabffab;
mem[2459] = 80'h0010ffabffabffabffab;
mem[2460] = 80'h0010ffabffabffabffab;
mem[2461] = 80'h0010ffabffabffabffab;
mem[2462] = 80'h0010ffabffabffabffab;
mem[2463] = 80'h0010ffabffabffabffab;
mem[2464] = 80'h0010ffabffabffabffab;
mem[2465] = 80'h0010ffabffabffabffab;
mem[2466] = 80'h0010ffabffabffabffab;
mem[2467] = 80'h0010ffabffabffabffab;
mem[2468] = 80'h0010ffabffabffabffab;
mem[2469] = 80'h0010ffabffabffabffab;
mem[2470] = 80'h0010ffabffabffabffab;
mem[2471] = 80'h0010ffabffabffabffab;
mem[2472] = 80'h0010ffabffabffabffab;
mem[2473] = 80'h0010ffabffabffabffab;
mem[2474] = 80'h0010ffabffabffabffab;
mem[2475] = 80'h0010ffabffabffabffab;
mem[2476] = 80'h0010ffabffabffabffab;
mem[2477] = 80'h0010ffabffabffabffab;
mem[2478] = 80'h0010ffabffabffabffab;
mem[2479] = 80'h0010ffabffabffabffab;
mem[2480] = 80'h0010ffabffabffabffab;
mem[2481] = 80'h0010ffabffabffabffab;
mem[2482] = 80'h0010ffabffabffabffab;
mem[2483] = 80'h0010ffabffabffabffab;
mem[2484] = 80'h0010ffabffabffabffab;
mem[2485] = 80'h0010ffabffabffabffab;
mem[2486] = 80'h0010ffabffabffabffab;
mem[2487] = 80'h0010ffabffabffabffab;
mem[2488] = 80'h0010ffabffabffabffab;
mem[2489] = 80'h0010ffabffabffabffab;
mem[2490] = 80'h0010ffabffabffabffab;
mem[2491] = 80'h0010ffabffabffabffab;
mem[2492] = 80'h0010ffabffabffabffab;
mem[2493] = 80'h0010ffabffabffabffab;
mem[2494] = 80'h0010ffabffabffabffab;
mem[2495] = 80'h0010ffabffabffabffab;
mem[2496] = 80'h0010ffabffabffabffab;
mem[2497] = 80'h0010ffabffabffabffab;
mem[2498] = 80'h0010ffabffabffabffab;
mem[2499] = 80'h0010ffabffabffabffab;
mem[2500] = 80'h0010ffabffabffabffab;
mem[2501] = 80'h0010ffabffabffabffab;
mem[2502] = 80'h0010ffabffabffabffab;
mem[2503] = 80'h0010ffabffabffabffab;
mem[2504] = 80'h0010ffabffabffabffab;
mem[2505] = 80'h0010ffabffabffabffab;
mem[2506] = 80'h0010ffabffabffabffab;
mem[2507] = 80'h0010ffabffabffabffab;
mem[2508] = 80'h0010ffabffabffabffab;
mem[2509] = 80'h0010ffabffabffabffab;
mem[2510] = 80'h0010ffabffabffabffab;
mem[2511] = 80'h0010ffabffabffabffab;
mem[2512] = 80'h0010ffabffabffabffab;
mem[2513] = 80'h0010ffabffabffabffab;
mem[2514] = 80'h0010ffabffabffabffab;
mem[2515] = 80'h0010ffabffabffabffab;
mem[2516] = 80'h0010ffabffabffabffab;
mem[2517] = 80'h0010ffabffabffabffab;
mem[2518] = 80'h0010ffabffabffabffab;
mem[2519] = 80'h0010ffabffabffabffab;
mem[2520] = 80'h0010ffabffabffabffab;
mem[2521] = 80'h0010ffabffabffabffab;
mem[2522] = 80'h0010ffabffabffabffab;
mem[2523] = 80'h0010ffabffabffabffab;
mem[2524] = 80'h0010ffabffabffabffab;
mem[2525] = 80'h0010ffabffabffabffab;
mem[2526] = 80'h0010ffabffabffabffab;
mem[2527] = 80'h0010ffabffabffabffab;
mem[2528] = 80'h0010ffabffabff4ead10;
mem[2529] = 80'h001048f8820687114a7f;
mem[2530] = 80'h0010d0126cbf5fbbc183;
mem[2531] = 80'h0115582ff7793a000000;
mem[2532] = 80'h10100000010000010010;
mem[2533] = 80'h00109400000208004500;
mem[2534] = 80'h0010015489b20000fffd;
mem[2535] = 80'h0010aea1c0550102c000;
mem[2536] = 80'h00100001ffabffabffab;
mem[2537] = 80'h0010ffabffabffabffab;
mem[2538] = 80'h0010ffabffabffabffab;
mem[2539] = 80'h0010ffabffabffabffab;
mem[2540] = 80'h0010ffabffabffabffab;
mem[2541] = 80'h0010ffabffabffabffab;
mem[2542] = 80'h0010ffabffabffabffab;
mem[2543] = 80'h0010ffabffabffabffab;
mem[2544] = 80'h0010ffabffabffabffab;
mem[2545] = 80'h0010ffabffabffabffab;
mem[2546] = 80'h0010ffabffabffabffab;
mem[2547] = 80'h0010ffabffabffabffab;
mem[2548] = 80'h0010ffabffabffabffab;
mem[2549] = 80'h0010ffabffabffabffab;
mem[2550] = 80'h0010ffabffabffabffab;
mem[2551] = 80'h0010ffabffabffabffab;
mem[2552] = 80'h0010ffabffabffabffab;
mem[2553] = 80'h0010ffabffabffabffab;
mem[2554] = 80'h0010ffabffabffabffab;
mem[2555] = 80'h0010ffabffabffabffab;
mem[2556] = 80'h0010ffabffabffabffab;
mem[2557] = 80'h0010ffabffabffabffab;
mem[2558] = 80'h0010ffabffabffabffab;
mem[2559] = 80'h0010ffabffabffabffab;
mem[2560] = 80'h0010ffabffabffabffab;
mem[2561] = 80'h0010ffabffabffabffab;
mem[2562] = 80'h0010ffabffabffabffab;
mem[2563] = 80'h0010ffabffabffabffab;
mem[2564] = 80'h0010ffabffabffabffab;
mem[2565] = 80'h0010ffabffabffabffab;
mem[2566] = 80'h0010ffabffabffabffab;
mem[2567] = 80'h0010ffabffabffabffab;
mem[2568] = 80'h0010ffabffabffabffab;
mem[2569] = 80'h0010ffabffabffabffab;
mem[2570] = 80'h0010ffabffabffabffab;
mem[2571] = 80'h0010ffabffabffabffab;
mem[2572] = 80'h0010ffabffabffabffab;
mem[2573] = 80'h0010ffabffabffab4d3f;
mem[2574] = 80'h0010723d900841474d3d;
mem[2575] = 80'h0010f7e60c1d39adbfb0;
mem[2576] = 80'h01162494281841e00000;
mem[2577] = 80'h10100000010000010010;
mem[2578] = 80'h00109400000208004500;
mem[2579] = 80'h001000bf89b30000fffd;
mem[2580] = 80'h0010af35c0550102c000;
mem[2581] = 80'h00100001ffabffabffab;
mem[2582] = 80'h0010ffabffabffabffab;
mem[2583] = 80'h0010ffabffabffabffab;
mem[2584] = 80'h0010ffabffabffabffab;
mem[2585] = 80'h0010ffabffabffabffab;
mem[2586] = 80'h0010ffabffabffabffab;
mem[2587] = 80'h0010ffabffabffabffab;
mem[2588] = 80'h0010ffabffabffabffab;
mem[2589] = 80'h0010ffabffabffabffab;
mem[2590] = 80'h0010ffabffabffabffab;
mem[2591] = 80'h0010ffabffabffabffab;
mem[2592] = 80'h0010ffabffabffabffab;
mem[2593] = 80'h0010ffabffabffabffab;
mem[2594] = 80'h0010ffabffabffabffab;
mem[2595] = 80'h0010ffabffabffabffab;
mem[2596] = 80'h0010ffabffabffabffab;
mem[2597] = 80'h0010ffabffabffabffab;
mem[2598] = 80'h0010ffabffabffabffab;
mem[2599] = 80'h0010ffabffabffabffab;
mem[2600] = 80'h0010ff4c4eac11487183;
mem[2601] = 80'h0010f886ef700bf9cd22;
mem[2602] = 80'h0010fc11f3157e2c1cf6;
mem[2603] = 80'h01111200000000000000;
mem[2604] = 80'h10100000010000010010;
mem[2605] = 80'h00109400000208004500;
mem[2606] = 80'h0010034c89b40000fffd;
mem[2607] = 80'h0010aca7c0550102c000;
mem[2608] = 80'h00100001ffabffabffab;
mem[2609] = 80'h0010ffabffabffabffab;
mem[2610] = 80'h0010ffabffabffabffab;
mem[2611] = 80'h0010ffabffabffabffab;
mem[2612] = 80'h0010ffabffabffabffab;
mem[2613] = 80'h0010ffabffabffabffab;
mem[2614] = 80'h0010ffabffabffabffab;
mem[2615] = 80'h0010ffabffabffabffab;
mem[2616] = 80'h0010ffabffabffabffab;
mem[2617] = 80'h0010ffabffabffabffab;
mem[2618] = 80'h0010ffabffabffabffab;
mem[2619] = 80'h0010ffabffabffabffab;
mem[2620] = 80'h0010ffabffabffabffab;
mem[2621] = 80'h0010ffabffabffabffab;
mem[2622] = 80'h0010ffabffabffabffab;
mem[2623] = 80'h0010ffabffabffabffab;
mem[2624] = 80'h0010ffabffabffabffab;
mem[2625] = 80'h0010ffabffabffabffab;
mem[2626] = 80'h0010ffabffabffabffab;
mem[2627] = 80'h0010ffabffabffabffab;
mem[2628] = 80'h0010ffabffabffabffab;
mem[2629] = 80'h0010ffabffabffabffab;
mem[2630] = 80'h0010ffabffabffabffab;
mem[2631] = 80'h0010ffabffabffabffab;
mem[2632] = 80'h0010ffabffabffabffab;
mem[2633] = 80'h0010ffabffabffabffab;
mem[2634] = 80'h0010ffabffabffabffab;
mem[2635] = 80'h0010ffabffabffabffab;
mem[2636] = 80'h0010ffabffabffabffab;
mem[2637] = 80'h0010ffabffabffabffab;
mem[2638] = 80'h0010ffabffabffabffab;
mem[2639] = 80'h0010ffabffabffabffab;
mem[2640] = 80'h0010ffabffabffabffab;
mem[2641] = 80'h0010ffabffabffabffab;
mem[2642] = 80'h0010ffabffabffabffab;
mem[2643] = 80'h0010ffabffabffabffab;
mem[2644] = 80'h0010ffabffabffabffab;
mem[2645] = 80'h0010ffabffabffabffab;
mem[2646] = 80'h0010ffabffabffabffab;
mem[2647] = 80'h0010ffabffabffabffab;
mem[2648] = 80'h0010ffabffabffabffab;
mem[2649] = 80'h0010ffabffabffabffab;
mem[2650] = 80'h0010ffabffabffabffab;
mem[2651] = 80'h0010ffabffabffabffab;
mem[2652] = 80'h0010ffabffabffabffab;
mem[2653] = 80'h0010ffabffabffabffab;
mem[2654] = 80'h0010ffabffabffabffab;
mem[2655] = 80'h0010ffabffabffabffab;
mem[2656] = 80'h0010ffabffabffabffab;
mem[2657] = 80'h0010ffabffabffabffab;
mem[2658] = 80'h0010ffabffabffabffab;
mem[2659] = 80'h0010ffabffabffabffab;
mem[2660] = 80'h0010ffabffabffabffab;
mem[2661] = 80'h0010ffabffabffabffab;
mem[2662] = 80'h0010ffabffabffabffab;
mem[2663] = 80'h0010ffabffabffabffab;
mem[2664] = 80'h0010ffabffabffabffab;
mem[2665] = 80'h0010ffabffabffabffab;
mem[2666] = 80'h0010ffabffabffabffab;
mem[2667] = 80'h0010ffabffabffabffab;
mem[2668] = 80'h0010ffabffabffabffab;
mem[2669] = 80'h0010ffabffabffabffab;
mem[2670] = 80'h0010ffabffabffabffab;
mem[2671] = 80'h0010ffabffabffabffab;
mem[2672] = 80'h0010ffabffabffabffab;
mem[2673] = 80'h0010ffabffabffabffab;
mem[2674] = 80'h0010ffabffabffabffab;
mem[2675] = 80'h0010ffabffabffabffab;
mem[2676] = 80'h0010ffabffabffabffab;
mem[2677] = 80'h0010ffabffabffabffab;
mem[2678] = 80'h0010ffabffabffabffab;
mem[2679] = 80'h0010ffabffabffabffab;
mem[2680] = 80'h0010ffabffabffabffab;
mem[2681] = 80'h0010ffabffabffabffab;
mem[2682] = 80'h0010ffabffabffabffab;
mem[2683] = 80'h0010ffabffabffabffab;
mem[2684] = 80'h0010ffabffabffabffab;
mem[2685] = 80'h0010ffabffabffabffab;
mem[2686] = 80'h0010ffabffabffabffab;
mem[2687] = 80'h0010ffabffabffabffab;
mem[2688] = 80'h0010ffabffabffabffab;
mem[2689] = 80'h0010ffabffabffabffab;
mem[2690] = 80'h0010ffabffabffabffab;
mem[2691] = 80'h0010ffabffabffabffab;
mem[2692] = 80'h0010ffabffabffabffab;
mem[2693] = 80'h0010ffabffabffabffab;
mem[2694] = 80'h0010ffabffabffabffab;
mem[2695] = 80'h0010ffabffabffabffab;
mem[2696] = 80'h0010ffabffabffabffab;
mem[2697] = 80'h0010ffabffabffabffab;
mem[2698] = 80'h0010ffabffabffabffab;
mem[2699] = 80'h0010ffabffabffabffab;
mem[2700] = 80'h0010ffabffabffabffab;
mem[2701] = 80'h0010ffabffabffabffab;
mem[2702] = 80'h0010ffabffabffabffab;
mem[2703] = 80'h0010ffabffabffabffab;
mem[2704] = 80'h0010ffabffabffabffab;
mem[2705] = 80'h0010ffabffabffabffab;
mem[2706] = 80'h0010ffabffabffabffab;
mem[2707] = 80'h0010ffabffabffabffab;
mem[2708] = 80'h0010ffabffabffab4b6a;
mem[2709] = 80'h001068fb99650c783e00;
mem[2710] = 80'h00106167c52cc61988da;
mem[2711] = 80'h0116f233cda47fee0000;
mem[2712] = 80'h10100000010000010010;
mem[2713] = 80'h00109400000208004500;
mem[2714] = 80'h001001bd89b50000fffd;
mem[2715] = 80'h0010ae35c0550102c000;
mem[2716] = 80'h00100001ffabffabffab;
mem[2717] = 80'h0010ffabffabffabffab;
mem[2718] = 80'h0010ffabffabffabffab;
mem[2719] = 80'h0010ffabffabffabffab;
mem[2720] = 80'h0010ffabffabffabffab;
mem[2721] = 80'h0010ffabffabffabffab;
mem[2722] = 80'h0010ffabffabffabffab;
mem[2723] = 80'h0010ffabffabffabffab;
mem[2724] = 80'h0010ffabffabffabffab;
mem[2725] = 80'h0010ffabffabffabffab;
mem[2726] = 80'h0010ffabffabffabffab;
mem[2727] = 80'h0010ffabffabffabffab;
mem[2728] = 80'h0010ffabffabffabffab;
mem[2729] = 80'h0010ffabffabffabffab;
mem[2730] = 80'h0010ffabffabffabffab;
mem[2731] = 80'h0010ffabffabffabffab;
mem[2732] = 80'h0010ffabffabffabffab;
mem[2733] = 80'h0010ffabffabffabffab;
mem[2734] = 80'h0010ffabffabffabffab;
mem[2735] = 80'h0010ffabffabffabffab;
mem[2736] = 80'h0010ffabffabffabffab;
mem[2737] = 80'h0010ffabffabffabffab;
mem[2738] = 80'h0010ffabffabffabffab;
mem[2739] = 80'h0010ffabffabffabffab;
mem[2740] = 80'h0010ffabffabffabffab;
mem[2741] = 80'h0010ffabffabffabffab;
mem[2742] = 80'h0010ffabffabffabffab;
mem[2743] = 80'h0010ffabffabffabffab;
mem[2744] = 80'h0010ffabffabffabffab;
mem[2745] = 80'h0010ffabffabffabffab;
mem[2746] = 80'h0010ffabffabffabffab;
mem[2747] = 80'h0010ffabffabffabffab;
mem[2748] = 80'h0010ffabffabffabffab;
mem[2749] = 80'h0010ffabffabffabffab;
mem[2750] = 80'h0010ffabffabffabffab;
mem[2751] = 80'h0010ffabffabffabffab;
mem[2752] = 80'h0010ffabffabffabffab;
mem[2753] = 80'h0010ffabffabffabffab;
mem[2754] = 80'h0010ffabffabffabffab;
mem[2755] = 80'h0010ffabffabffabffab;
mem[2756] = 80'h0010ffabffabffabffab;
mem[2757] = 80'h0010ffabffabffabffab;
mem[2758] = 80'h0010ffabffabffabffab;
mem[2759] = 80'h0010ffabffabffabffab;
mem[2760] = 80'h0010ffabffabffabffab;
mem[2761] = 80'h0010ffabffabffabffab;
mem[2762] = 80'h0010ffabffabffabffab;
mem[2763] = 80'h0010ffabffabffabffab;
mem[2764] = 80'h0010ffabffabffabffab;
mem[2765] = 80'h0010ffabffabffabffab;
mem[2766] = 80'h0010ffabffabffabff4a;
mem[2767] = 80'h00101bb6d7411ccec7f5;
mem[2768] = 80'h0010d2e68a30fb854824;
mem[2769] = 80'h01171f386818eabdf300;
mem[2770] = 80'h10100000010000010010;
mem[2771] = 80'h00109400000208004500;
mem[2772] = 80'h001000f589b60000fffd;
mem[2773] = 80'h0010aefcc0550102c000;
mem[2774] = 80'h00100001ffabffabffab;
mem[2775] = 80'h0010ffabffabffabffab;
mem[2776] = 80'h0010ffabffabffabffab;
mem[2777] = 80'h0010ffabffabffabffab;
mem[2778] = 80'h0010ffabffabffabffab;
mem[2779] = 80'h0010ffabffabffabffab;
mem[2780] = 80'h0010ffabffabffabffab;
mem[2781] = 80'h0010ffabffabffabffab;
mem[2782] = 80'h0010ffabffabffabffab;
mem[2783] = 80'h0010ffabffabffabffab;
mem[2784] = 80'h0010ffabffabffabffab;
mem[2785] = 80'h0010ffabffabffabffab;
mem[2786] = 80'h0010ffabffabffabffab;
mem[2787] = 80'h0010ffabffabffabffab;
mem[2788] = 80'h0010ffabffabffabffab;
mem[2789] = 80'h0010ffabffabffabffab;
mem[2790] = 80'h0010ffabffabffabffab;
mem[2791] = 80'h0010ffabffabffabffab;
mem[2792] = 80'h0010ffabffabffabffab;
mem[2793] = 80'h0010ffabffabffabffab;
mem[2794] = 80'h0010ffabffabffabffab;
mem[2795] = 80'h0010ffabffabffabffab;
mem[2796] = 80'h0010ffabffabffabffab;
mem[2797] = 80'h0010ffabffabffabffab;
mem[2798] = 80'h0010ffabffabffabffab;
mem[2799] = 80'h0010ffabffabffabff49;
mem[2800] = 80'h001089d4a229968907a9;
mem[2801] = 80'h0010a56ebc2e8ab7baf2;
mem[2802] = 80'h0117a73de7c4a4349e00;
mem[2803] = 80'h10100000010000010010;
mem[2804] = 80'h00109400000208004500;
mem[2805] = 80'h0010036a89b70000fffd;
mem[2806] = 80'h0010ac86c0550102c000;
mem[2807] = 80'h00100001ffabffabffab;
mem[2808] = 80'h0010ffabffabffabffab;
mem[2809] = 80'h0010ffabffabffabffab;
mem[2810] = 80'h0010ffabffabffabffab;
mem[2811] = 80'h0010ffabffabffabffab;
mem[2812] = 80'h0010ffabffabffabffab;
mem[2813] = 80'h0010ffabffabffabffab;
mem[2814] = 80'h0010ffabffabffabffab;
mem[2815] = 80'h0010ffabffabffabffab;
mem[2816] = 80'h0010ffabffabffabffab;
mem[2817] = 80'h0010ffabffabffabffab;
mem[2818] = 80'h0010ffabffabffabffab;
mem[2819] = 80'h0010ffabffabffabffab;
mem[2820] = 80'h0010ffabffabffabffab;
mem[2821] = 80'h0010ffabffabffabffab;
mem[2822] = 80'h0010ffabffabffabffab;
mem[2823] = 80'h0010ffabffabffabffab;
mem[2824] = 80'h0010ffabffabffabffab;
mem[2825] = 80'h0010ffabffabffabffab;
mem[2826] = 80'h0010ffabffabffabffab;
mem[2827] = 80'h0010ffabffabffabffab;
mem[2828] = 80'h0010ffabffabffabffab;
mem[2829] = 80'h0010ffabffabffabffab;
mem[2830] = 80'h0010ffabffabffabffab;
mem[2831] = 80'h0010ffabffabffabffab;
mem[2832] = 80'h0010ffabffabffabffab;
mem[2833] = 80'h0010ffabffabffabffab;
mem[2834] = 80'h0010ffabffabffabffab;
mem[2835] = 80'h0010ffabffabffabffab;
mem[2836] = 80'h0010ffabffabffabffab;
mem[2837] = 80'h0010ffabffabffabffab;
mem[2838] = 80'h0010ffabffabffabffab;
mem[2839] = 80'h0010ffabffabffabffab;
mem[2840] = 80'h0010ffabffabffabffab;
mem[2841] = 80'h0010ffabffabffabffab;
mem[2842] = 80'h0010ffabffabffabffab;
mem[2843] = 80'h0010ffabffabffabffab;
mem[2844] = 80'h0010ffabffabffabffab;
mem[2845] = 80'h0010ffabffabffabffab;
mem[2846] = 80'h0010ffabffabffabffab;
mem[2847] = 80'h0010ffabffabffabffab;
mem[2848] = 80'h0010ffabffabffabffab;
mem[2849] = 80'h0010ffabffabffabffab;
mem[2850] = 80'h0010ffabffabffabffab;
mem[2851] = 80'h0010ffabffabffabffab;
mem[2852] = 80'h0010ffabffabffabffab;
mem[2853] = 80'h0010ffabffabffabffab;
mem[2854] = 80'h0010ffabffabffabffab;
mem[2855] = 80'h0010ffabffabffabffab;
mem[2856] = 80'h0010ffabffabffabffab;
mem[2857] = 80'h0010ffabffabffabffab;
mem[2858] = 80'h0010ffabffabffabffab;
mem[2859] = 80'h0010ffabffabffabffab;
mem[2860] = 80'h0010ffabffabffabffab;
mem[2861] = 80'h0010ffabffabffabffab;
mem[2862] = 80'h0010ffabffabffabffab;
mem[2863] = 80'h0010ffabffabffabffab;
mem[2864] = 80'h0010ffabffabffabffab;
mem[2865] = 80'h0010ffabffabffabffab;
mem[2866] = 80'h0010ffabffabffabffab;
mem[2867] = 80'h0010ffabffabffabffab;
mem[2868] = 80'h0010ffabffabffabffab;
mem[2869] = 80'h0010ffabffabffabffab;
mem[2870] = 80'h0010ffabffabffabffab;
mem[2871] = 80'h0010ffabffabffabffab;
mem[2872] = 80'h0010ffabffabffabffab;
mem[2873] = 80'h0010ffabffabffabffab;
mem[2874] = 80'h0010ffabffabffabffab;
mem[2875] = 80'h0010ffabffabffabffab;
mem[2876] = 80'h0010ffabffabffabffab;
mem[2877] = 80'h0010ffabffabffabffab;
mem[2878] = 80'h0010ffabffabffabffab;
mem[2879] = 80'h0010ffabffabffabffab;
mem[2880] = 80'h0010ffabffabffabffab;
mem[2881] = 80'h0010ffabffabffabffab;
mem[2882] = 80'h0010ffabffabffabffab;
mem[2883] = 80'h0010ffabffabffabffab;
mem[2884] = 80'h0010ffabffabffabffab;
mem[2885] = 80'h0010ffabffabffabffab;
mem[2886] = 80'h0010ffabffabffabffab;
mem[2887] = 80'h0010ffabffabffabffab;
mem[2888] = 80'h0010ffabffabffabffab;
mem[2889] = 80'h0010ffabffabffabffab;
mem[2890] = 80'h0010ffabffabffabffab;
mem[2891] = 80'h0010ffabffabffabffab;
mem[2892] = 80'h0010ffabffabffabffab;
mem[2893] = 80'h0010ffabffabffabffab;
mem[2894] = 80'h0010ffabffabffabffab;
mem[2895] = 80'h0010ffabffabffabffab;
mem[2896] = 80'h0010ffabffabffabffab;
mem[2897] = 80'h0010ffabffabffabffab;
mem[2898] = 80'h0010ffabffabffabffab;
mem[2899] = 80'h0010ffabffabffabffab;
mem[2900] = 80'h0010ffabffabffabffab;
mem[2901] = 80'h0010ffabffabffabffab;
mem[2902] = 80'h0010ffabffabffabffab;
mem[2903] = 80'h0010ffabffabffabffab;
mem[2904] = 80'h0010ffabffabffabffab;
mem[2905] = 80'h0010ffabffabffabffab;
mem[2906] = 80'h0010ffabffabffabffab;
mem[2907] = 80'h0010ffabffabffabffab;
mem[2908] = 80'h0010ffabffabffabffab;
mem[2909] = 80'h0010ffabffabffabffab;
mem[2910] = 80'h0010ffabffabffabffab;
mem[2911] = 80'h0010ffabffab48f80a8e;
mem[2912] = 80'h0010f1ef4bb86277e951;
mem[2913] = 80'h0010db5a79ebb636178b;
mem[2914] = 80'h01140fb7e9bb00000000;
mem[2915] = 80'h10100000010000010010;
mem[2916] = 80'h00109400000208004500;
mem[2917] = 80'h001004a289b80000fffd;
mem[2918] = 80'h0010ab4dc0550102c000;
mem[2919] = 80'h00100001ffabffabffab;
mem[2920] = 80'h0010ffabffabffabffab;
mem[2921] = 80'h0010ffabffabffabffab;
mem[2922] = 80'h0010ffabffabffabffab;
mem[2923] = 80'h0010ffabffabffabffab;
mem[2924] = 80'h0010ffabffabffabffab;
mem[2925] = 80'h0010ffabffabffabffab;
mem[2926] = 80'h0010ffabffabffabffab;
mem[2927] = 80'h0010ffabffabffabffab;
mem[2928] = 80'h0010ffabffabffabffab;
mem[2929] = 80'h0010ffabffabffabffab;
mem[2930] = 80'h0010ffabffabffabffab;
mem[2931] = 80'h0010ffabffabffabffab;
mem[2932] = 80'h0010ffabffabffabffab;
mem[2933] = 80'h0010ffabffabffabffab;
mem[2934] = 80'h0010ffabffabffabffab;
mem[2935] = 80'h0010ffabffabffabffab;
mem[2936] = 80'h0010ffabffabffabffab;
mem[2937] = 80'h0010ffabffabffabffab;
mem[2938] = 80'h0010ffabffabffabffab;
mem[2939] = 80'h0010ffabffabffabffab;
mem[2940] = 80'h0010ffabffabffabffab;
mem[2941] = 80'h0010ffabffabffabffab;
mem[2942] = 80'h0010ffabffabffabffab;
mem[2943] = 80'h0010ffabffabffabffab;
mem[2944] = 80'h0010ffabffabffabffab;
mem[2945] = 80'h0010ffabffabffabffab;
mem[2946] = 80'h0010ffabffabffabffab;
mem[2947] = 80'h0010ffabffabffabffab;
mem[2948] = 80'h0010ffabffabffabffab;
mem[2949] = 80'h0010ffabffabffabffab;
mem[2950] = 80'h0010ffabffabffabffab;
mem[2951] = 80'h0010ffabffabffabffab;
mem[2952] = 80'h0010ffabffabffabffab;
mem[2953] = 80'h0010ffabffabffabffab;
mem[2954] = 80'h0010ffabffabffabffab;
mem[2955] = 80'h0010ffabffabffabffab;
mem[2956] = 80'h0010ffabffabffabffab;
mem[2957] = 80'h0010ffabffabffabffab;
mem[2958] = 80'h0010ffabffabffabffab;
mem[2959] = 80'h0010ffabffabffabffab;
mem[2960] = 80'h0010ffabffabffabffab;
mem[2961] = 80'h0010ffabffabffabffab;
mem[2962] = 80'h0010ffabffabffabffab;
mem[2963] = 80'h0010ffabffabffabffab;
mem[2964] = 80'h0010ffabffabffabffab;
mem[2965] = 80'h0010ffabffabffabffab;
mem[2966] = 80'h0010ffabffabffabffab;
mem[2967] = 80'h0010ffabffabffabffab;
mem[2968] = 80'h0010ffabffabffabffab;
mem[2969] = 80'h0010ffabffabffabffab;
mem[2970] = 80'h0010ffabffabffabffab;
mem[2971] = 80'h0010ffabffabffabffab;
mem[2972] = 80'h0010ffabffabffabffab;
mem[2973] = 80'h0010ffabffabffabffab;
mem[2974] = 80'h0010ffabffabffabffab;
mem[2975] = 80'h0010ffabffabffabffab;
mem[2976] = 80'h0010ffabffabffabffab;
mem[2977] = 80'h0010ffabffabffabffab;
mem[2978] = 80'h0010ffabffabffabffab;
mem[2979] = 80'h0010ffabffabffabffab;
mem[2980] = 80'h0010ffabffabffabffab;
mem[2981] = 80'h0010ffabffabffabffab;
mem[2982] = 80'h0010ffabffabffabffab;
mem[2983] = 80'h0010ffabffabffabffab;
mem[2984] = 80'h0010ffabffabffabffab;
mem[2985] = 80'h0010ffabffabffabffab;
mem[2986] = 80'h0010ffabffabffabffab;
mem[2987] = 80'h0010ffabffabffabffab;
mem[2988] = 80'h0010ffabffabffabffab;
mem[2989] = 80'h0010ffabffabffabffab;
mem[2990] = 80'h0010ffabffabffabffab;
mem[2991] = 80'h0010ffabffabffabffab;
mem[2992] = 80'h0010ffabffabffabffab;
mem[2993] = 80'h0010ffabffabffabffab;
mem[2994] = 80'h0010ffabffabffabffab;
mem[2995] = 80'h0010ffabffabffabffab;
mem[2996] = 80'h0010ffabffabffabffab;
mem[2997] = 80'h0010ffabffabffabffab;
mem[2998] = 80'h0010ffabffabffabffab;
mem[2999] = 80'h0010ffabffabffabffab;
mem[3000] = 80'h0010ffabffabffabffab;
mem[3001] = 80'h0010ffabffabffabffab;
mem[3002] = 80'h0010ffabffabffabffab;
mem[3003] = 80'h0010ffabffabffabffab;
mem[3004] = 80'h0010ffabffabffabffab;
mem[3005] = 80'h0010ffabffabffabffab;
mem[3006] = 80'h0010ffabffabffabffab;
mem[3007] = 80'h0010ffabffabffabffab;
mem[3008] = 80'h0010ffabffabffabffab;
mem[3009] = 80'h0010ffabffabffabffab;
mem[3010] = 80'h0010ffabffabffabffab;
mem[3011] = 80'h0010ffabffabffabffab;
mem[3012] = 80'h0010ffabffabffabffab;
mem[3013] = 80'h0010ffabffabffabffab;
mem[3014] = 80'h0010ffabffabffabffab;
mem[3015] = 80'h0010ffabffabffabffab;
mem[3016] = 80'h0010ffabffabffabffab;
mem[3017] = 80'h0010ffabffabffabffab;
mem[3018] = 80'h0010ffabffabffabffab;
mem[3019] = 80'h0010ffabffabffabffab;
mem[3020] = 80'h0010ffabffabffabffab;
mem[3021] = 80'h0010ffabffabffabffab;
mem[3022] = 80'h0010ffabffabffabffab;
mem[3023] = 80'h0010ffabffabffabffab;
mem[3024] = 80'h0010ffabffabffabffab;
mem[3025] = 80'h0010ffabffabffabffab;
mem[3026] = 80'h0010ffabffabffabffab;
mem[3027] = 80'h0010ffabffabffabffab;
mem[3028] = 80'h0010ffabffabffabffab;
mem[3029] = 80'h0010ffabffabffabffab;
mem[3030] = 80'h0010ffabffabffabffab;
mem[3031] = 80'h0010ffabffabffabffab;
mem[3032] = 80'h0010ffabffabffabffab;
mem[3033] = 80'h0010ffabffabffabffab;
mem[3034] = 80'h0010ffabffabffabffab;
mem[3035] = 80'h0010ffabffabffabffab;
mem[3036] = 80'h0010ffabffabffabffab;
mem[3037] = 80'h0010ffabffabffabffab;
mem[3038] = 80'h0010ffabffabffabffab;
mem[3039] = 80'h0010ffabffabffabffab;
mem[3040] = 80'h0010ffabffabffabffab;
mem[3041] = 80'h0010ffabffabffabffab;
mem[3042] = 80'h0010ffabffabffabffab;
mem[3043] = 80'h0010ffabffabffabffab;
mem[3044] = 80'h0010ffabffabffabffab;
mem[3045] = 80'h0010ffabffabffabffab;
mem[3046] = 80'h0010ffabffabffabffab;
mem[3047] = 80'h0010ffabffabffabffab;
mem[3048] = 80'h0010ffabffabffabffab;
mem[3049] = 80'h0010ffabffabffabffab;
mem[3050] = 80'h0010ffabffabffabffab;
mem[3051] = 80'h0010ffabffabffabffab;
mem[3052] = 80'h0010ffabffabffabffab;
mem[3053] = 80'h0010ffabffabffabffab;
mem[3054] = 80'h0010ffabffabffabffab;
mem[3055] = 80'h0010ffabffabffabffab;
mem[3056] = 80'h0010ffabffabffabffab;
mem[3057] = 80'h0010ffabffabffabffab;
mem[3058] = 80'h0010ffabffabffabffab;
mem[3059] = 80'h0010ffabffabffabffab;
mem[3060] = 80'h0010ffabffabffabffab;
mem[3061] = 80'h0010ffabffabffabffab;
mem[3062] = 80'h0010ffabffab47c05d77;
mem[3063] = 80'h00108bbf9606d87b4c64;
mem[3064] = 80'h0010574b887117f21c73;
mem[3065] = 80'h01148bc002c700000000;
mem[3066] = 80'h00000000000000000000;
mem[3067] = 80'h00000000000000000000;
mem[3068] = 80'h00000000000000000000;
mem[3069] = 80'h00000000000000000000;
mem[3070] = 80'h00000000000000000000;
mem[3071] = 80'h00000000000000000000;
mem[3072] = 80'h00000000000000000000;
mem[3073] = 80'h00000000000000000000;
mem[3074] = 80'h00000000000000000000;
mem[3075] = 80'h00000000000000000000;
mem[3076] = 80'h00000000000000000000;
mem[3077] = 80'h00000000000000000000;
mem[3078] = 80'h00000000000000000000;
mem[3079] = 80'h00000000000000000000;
mem[3080] = 80'h00000000000000000000;
mem[3081] = 80'h00000000000000000000;
mem[3082] = 80'h10100000010000010010;
mem[3083] = 80'h00109400000208004500;
mem[3084] = 80'h0010053e89b90000fffd;
mem[3085] = 80'h0010aab0c0550102c000;
mem[3086] = 80'h00100001ffabffabffab;
mem[3087] = 80'h0010ffabffabffabffab;
mem[3088] = 80'h0010ffabffabffabffab;
mem[3089] = 80'h0010ffabffabffabffab;
mem[3090] = 80'h0010ffabffabffabffab;
mem[3091] = 80'h0010ffabffabffabffab;
mem[3092] = 80'h0010ffabffabffabffab;
mem[3093] = 80'h0010ffabffabffabffab;
mem[3094] = 80'h0010ffabffabffabffab;
mem[3095] = 80'h0010ffabffabffabffab;
mem[3096] = 80'h0010ffabffabffabffab;
mem[3097] = 80'h0010ffabffabffabffab;
mem[3098] = 80'h0010ffabffabffabffab;
mem[3099] = 80'h0010ffabffabffabffab;
mem[3100] = 80'h0010ffabffabffabffab;
mem[3101] = 80'h0010ffabffabffabffab;
mem[3102] = 80'h0010ffabffabffabffab;
mem[3103] = 80'h0010ffabffabffabffab;
mem[3104] = 80'h0010ffabffabffabffab;
mem[3105] = 80'h0010ffabffabffabffab;
mem[3106] = 80'h0010ffabffabffabffab;
mem[3107] = 80'h0010ffabffabffabffab;
mem[3108] = 80'h0010ffabffabffabffab;
mem[3109] = 80'h0010ffabffabffabffab;
mem[3110] = 80'h0010ffabffabffabffab;
mem[3111] = 80'h0010ffabffabffabffab;
mem[3112] = 80'h0010ffabffabffabffab;
mem[3113] = 80'h0010ffabffabffabffab;
mem[3114] = 80'h0010ffabffabffabffab;
mem[3115] = 80'h0010ffabffabffabffab;
mem[3116] = 80'h0010ffabffabffabffab;
mem[3117] = 80'h0010ffabffabffabffab;
mem[3118] = 80'h0010ffabffabffabffab;
mem[3119] = 80'h0010ffabffabffabffab;
mem[3120] = 80'h0010ffabffabffabffab;
mem[3121] = 80'h0010ffabffabffabffab;
mem[3122] = 80'h0010ffabffabffabffab;
mem[3123] = 80'h0010ffabffabffabffab;
mem[3124] = 80'h0010ffabffabffabffab;
mem[3125] = 80'h0010ffabffabffabffab;
mem[3126] = 80'h0010ffabffabffabffab;
mem[3127] = 80'h0010ffabffabffabffab;
mem[3128] = 80'h0010ffabffabffabffab;
mem[3129] = 80'h0010ffabffabffabffab;
mem[3130] = 80'h0010ffabffabffabffab;
mem[3131] = 80'h0010ffabffabffabffab;
mem[3132] = 80'h0010ffabffabffabffab;
mem[3133] = 80'h0010ffabffabffabffab;
mem[3134] = 80'h0010ffabffabffabffab;
mem[3135] = 80'h0010ffabffabffabffab;
mem[3136] = 80'h0010ffabffabffabffab;
mem[3137] = 80'h0010ffabffabffabffab;
mem[3138] = 80'h0010ffabffabffabffab;
mem[3139] = 80'h0010ffabffabffabffab;
mem[3140] = 80'h0010ffabffabffabffab;
mem[3141] = 80'h0010ffabffabffabffab;
mem[3142] = 80'h0010ffabffabffabffab;
mem[3143] = 80'h0010ffabffabffabffab;
mem[3144] = 80'h0010ffabffabffabffab;
mem[3145] = 80'h0010ffabffabffabffab;
mem[3146] = 80'h0010ffabffabffabffab;
mem[3147] = 80'h0010ffabffabffabffab;
mem[3148] = 80'h0010ffabffabffabffab;
mem[3149] = 80'h0010ffabffabffabffab;
mem[3150] = 80'h0010ffabffabffabffab;
mem[3151] = 80'h0010ffabffabffabffab;
mem[3152] = 80'h0010ffabffabffabffab;
mem[3153] = 80'h0010ffabffabffabffab;
mem[3154] = 80'h0010ffabffabffabffab;
mem[3155] = 80'h0010ffabffabffabffab;
mem[3156] = 80'h0010ffabffabffabffab;
mem[3157] = 80'h0010ffabffabffabffab;
mem[3158] = 80'h0010ffabffabffabffab;
mem[3159] = 80'h0010ffabffabffabffab;
mem[3160] = 80'h0010ffabffabffabffab;
mem[3161] = 80'h0010ffabffabffabffab;
mem[3162] = 80'h0010ffabffabffabffab;
mem[3163] = 80'h0010ffabffabffabffab;
mem[3164] = 80'h0010ffabffabffabffab;
mem[3165] = 80'h0010ffabffabffabffab;
mem[3166] = 80'h0010ffabffabffabffab;
mem[3167] = 80'h0010ffabffabffabffab;
mem[3168] = 80'h0010ffabffabffabffab;
mem[3169] = 80'h0010ffabffabffabffab;
mem[3170] = 80'h0010ffabffabffabffab;
mem[3171] = 80'h0010ffabffabffabffab;
mem[3172] = 80'h0010ffabffabffabffab;
mem[3173] = 80'h0010ffabffabffabffab;
mem[3174] = 80'h0010ffabffabffabffab;
mem[3175] = 80'h0010ffabffabffabffab;
mem[3176] = 80'h0010ffabffabffabffab;
mem[3177] = 80'h0010ffabffabffabffab;
mem[3178] = 80'h0010ffabffabffabffab;
mem[3179] = 80'h0010ffabffabffabffab;
mem[3180] = 80'h0010ffabffabffabffab;
mem[3181] = 80'h0010ffabffabffabffab;
mem[3182] = 80'h0010ffabffabffabffab;
mem[3183] = 80'h0010ffabffabffabffab;
mem[3184] = 80'h0010ffabffabffabffab;
mem[3185] = 80'h0010ffabffabffabffab;
mem[3186] = 80'h0010ffabffabffabffab;
mem[3187] = 80'h0010ffabffabffabffab;
mem[3188] = 80'h0010ffabffabffabffab;
mem[3189] = 80'h0010ffabffabffabffab;
mem[3190] = 80'h0010ffabffabffabffab;
mem[3191] = 80'h0010ffabffabffabffab;
mem[3192] = 80'h0010ffabffabffabffab;
mem[3193] = 80'h0010ffabffabffabffab;
mem[3194] = 80'h0010ffabffabffabffab;
mem[3195] = 80'h0010ffabffabffabffab;
mem[3196] = 80'h0010ffabffabffabffab;
mem[3197] = 80'h0010ffabffabffabffab;
mem[3198] = 80'h0010ffabffabffabffab;
mem[3199] = 80'h0010ffabffabffabffab;
mem[3200] = 80'h0010ffabffabffabffab;
mem[3201] = 80'h0010ffabffabffabffab;
mem[3202] = 80'h0010ffabffabffabffab;
mem[3203] = 80'h0010ffabffabffabffab;
mem[3204] = 80'h0010ffabffabffabffab;
mem[3205] = 80'h0010ffabffabffabffab;
mem[3206] = 80'h0010ffabffabffabffab;
mem[3207] = 80'h0010ffabffabffabffab;
mem[3208] = 80'h0010ffabffabffabffab;
mem[3209] = 80'h0010ffabffabffabffab;
mem[3210] = 80'h0010ffabffabffabffab;
mem[3211] = 80'h0010ffabffabffabffab;
mem[3212] = 80'h0010ffabffabffabffab;
mem[3213] = 80'h0010ffabffabffabffab;
mem[3214] = 80'h0010ffabffabffabffab;
mem[3215] = 80'h0010ffabffabffabffab;
mem[3216] = 80'h0010ffabffabffabffab;
mem[3217] = 80'h0010ffabffabffabffab;
mem[3218] = 80'h0010ffabffabffabffab;
mem[3219] = 80'h0010ffabffabffabffab;
mem[3220] = 80'h0010ffabffabffabffab;
mem[3221] = 80'h0010ffabffabffabffab;
mem[3222] = 80'h0010ffabffabffabffab;
mem[3223] = 80'h0010ffabffabffabffab;
mem[3224] = 80'h0010ffabffabffabffab;
mem[3225] = 80'h0010ffabffabffabffab;
mem[3226] = 80'h0010ffabffabffabffab;
mem[3227] = 80'h0010ffabffabffabffab;
mem[3228] = 80'h0010ffabffabffabffab;
mem[3229] = 80'h0010ffabffabffabffab;
mem[3230] = 80'h0010ffabffabffabffab;
mem[3231] = 80'h0010ffabffabffabffab;
mem[3232] = 80'h0010ffabffabffabffab;
mem[3233] = 80'h0010ffabffabffabffab;
mem[3234] = 80'h0010ffabffabffabffab;
mem[3235] = 80'h0010ffabffabffabffab;
mem[3236] = 80'h0010ffabffabffabffab;
mem[3237] = 80'h0010ffabffabffabffab;
mem[3238] = 80'h0010ffabffabffabffab;
mem[3239] = 80'h0010ffabffabffabffab;
mem[3240] = 80'h0010ffabffabffabffab;
mem[3241] = 80'h0010ffabffabffabffab;
mem[3242] = 80'h0010ffabffabffabffab;
mem[3243] = 80'h0010ffabffabffabffab;
mem[3244] = 80'h0010ffabffabffabffab;
mem[3245] = 80'h0010ffabffabffabffab;
mem[3246] = 80'h0010ffabffabffabffab;
mem[3247] = 80'h0010ffabffabffabffab;
mem[3248] = 80'h0010ffabffabffabffab;
mem[3249] = 80'h001046b1835b53c654b9;
mem[3250] = 80'h001013a9cb89a2959420;
mem[3251] = 80'h01103b273c63d547be4f;
mem[3252] = 80'h10100000010000010010;
mem[3253] = 80'h00109400000208004500;
mem[3254] = 80'h001002b689ba0000fffd;
mem[3255] = 80'h0010ad37c0550102c000;
mem[3256] = 80'h00100001ffabffabffab;
mem[3257] = 80'h0010ffabffabffabffab;
mem[3258] = 80'h0010ffabffabffabffab;
mem[3259] = 80'h0010ffabffabffabffab;
mem[3260] = 80'h0010ffabffabffabffab;
mem[3261] = 80'h0010ffabffabffabffab;
mem[3262] = 80'h0010ffabffabffabffab;
mem[3263] = 80'h0010ffabffabffabffab;
mem[3264] = 80'h0010ffabffabffabffab;
mem[3265] = 80'h0010ffabffabffabffab;
mem[3266] = 80'h0010ffabffabffabffab;
mem[3267] = 80'h0010ffabffabffabffab;
mem[3268] = 80'h0010ffabffabffabffab;
mem[3269] = 80'h0010ffabffabffabffab;
mem[3270] = 80'h0010ffabffabffabffab;
mem[3271] = 80'h0010ffabffabffabffab;
mem[3272] = 80'h0010ffabffabffabffab;
mem[3273] = 80'h0010ffabffabffabffab;
mem[3274] = 80'h0010ffabffabffabffab;
mem[3275] = 80'h0010ffabffabffabffab;
mem[3276] = 80'h0010ffabffabffabffab;
mem[3277] = 80'h0010ffabffabffabffab;
mem[3278] = 80'h0010ffabffabffabffab;
mem[3279] = 80'h0010ffabffabffabffab;
mem[3280] = 80'h0010ffabffabffabffab;
mem[3281] = 80'h0010ffabffabffabffab;
mem[3282] = 80'h0010ffabffabffabffab;
mem[3283] = 80'h0010ffabffabffabffab;
mem[3284] = 80'h0010ffabffabffabffab;
mem[3285] = 80'h0010ffabffabffabffab;
mem[3286] = 80'h0010ffabffabffabffab;
mem[3287] = 80'h0010ffabffabffabffab;
mem[3288] = 80'h0010ffabffabffabffab;
mem[3289] = 80'h0010ffabffabffabffab;
mem[3290] = 80'h0010ffabffabffabffab;
mem[3291] = 80'h0010ffabffabffabffab;
mem[3292] = 80'h0010ffabffabffabffab;
mem[3293] = 80'h0010ffabffabffabffab;
mem[3294] = 80'h0010ffabffabffabffab;
mem[3295] = 80'h0010ffabffabffabffab;
mem[3296] = 80'h0010ffabffabffabffab;
mem[3297] = 80'h0010ffabffabffabffab;
mem[3298] = 80'h0010ffabffabffabffab;
mem[3299] = 80'h0010ffabffabffabffab;
mem[3300] = 80'h0010ffabffabffabffab;
mem[3301] = 80'h0010ffabffabffabffab;
mem[3302] = 80'h0010ffabffabffabffab;
mem[3303] = 80'h0010ffabffabffabffab;
mem[3304] = 80'h0010ffabffabffabffab;
mem[3305] = 80'h0010ffabffabffabffab;
mem[3306] = 80'h0010ffabffabffabffab;
mem[3307] = 80'h0010ffabffabffabffab;
mem[3308] = 80'h0010ffabffabffabffab;
mem[3309] = 80'h0010ffabffabffabffab;
mem[3310] = 80'h0010ffabffabffabffab;
mem[3311] = 80'h0010ffabffabffabffab;
mem[3312] = 80'h0010ffabffabffabffab;
mem[3313] = 80'h0010ffabffabffabffab;
mem[3314] = 80'h0010ffabffabffabffab;
mem[3315] = 80'h0010ffabffabffabffab;
mem[3316] = 80'h0010ffabffabffabffab;
mem[3317] = 80'h0010ffabffabffabffab;
mem[3318] = 80'h0010ffabffabffabffab;
mem[3319] = 80'h0010ffabffabffabffab;
mem[3320] = 80'h0010ffabffabffabffab;
mem[3321] = 80'h0010ffabffabffabffab;
mem[3322] = 80'h0010ffabffabffabffab;
mem[3323] = 80'h0010ffabffabffabffab;
mem[3324] = 80'h0010ffabffabffabffab;
mem[3325] = 80'h0010ffabffabffabffab;
mem[3326] = 80'h0010ffabffabffabffab;
mem[3327] = 80'h0010ffabffabffabffab;
mem[3328] = 80'h0010ffabffabffabffab;
mem[3329] = 80'h0010ffabffabffabffab;
mem[3330] = 80'h0010ffabffabffabffab;
mem[3331] = 80'h0010ffabffabffabffab;
mem[3332] = 80'h0010ffabffabffabffab;
mem[3333] = 80'h0010ffabffabffabffab;
mem[3334] = 80'h0010ffabffabffabffab;
mem[3335] = 80'h0010ffabffabffabffab;
mem[3336] = 80'h0010ffabffabffabffab;
mem[3337] = 80'h0010ffabffabffabffab;
mem[3338] = 80'h00104523e12e3b4c1379;
mem[3339] = 80'h00104fde43bfbce7fed2;
mem[3340] = 80'h011033d907b72f689772;
mem[3341] = 80'h10100000010000010010;
mem[3342] = 80'h00109400000208004500;
mem[3343] = 80'h0010044b89bb0000fffd;
mem[3344] = 80'h0010aba1c0550102c000;
mem[3345] = 80'h00100001ffabffabffab;
mem[3346] = 80'h0010ffabffabffabffab;
mem[3347] = 80'h0010ffabffabffabffab;
mem[3348] = 80'h0010ffabffabffabffab;
mem[3349] = 80'h0010ffabffabffabffab;
mem[3350] = 80'h0010ffabffabffabffab;
mem[3351] = 80'h0010ffabffabffabffab;
mem[3352] = 80'h0010ffabffabffabffab;
mem[3353] = 80'h0010ffabffabffabffab;
mem[3354] = 80'h0010ffabffabffabffab;
mem[3355] = 80'h0010ffabffabffabffab;
mem[3356] = 80'h0010ffabffabffabffab;
mem[3357] = 80'h0010ffabffabffabffab;
mem[3358] = 80'h0010ffabffabffabffab;
mem[3359] = 80'h0010ffabffabffabffab;
mem[3360] = 80'h0010ffabffabffabffab;
mem[3361] = 80'h0010ffabffabffabffab;
mem[3362] = 80'h0010ffabffabffabffab;
mem[3363] = 80'h0010ffabffabffabffab;
mem[3364] = 80'h0010ffabffabffabffab;
mem[3365] = 80'h0010ffabffabffabffab;
mem[3366] = 80'h0010ffabffabffabffab;
mem[3367] = 80'h0010ffabffabffabffab;
mem[3368] = 80'h0010ffabffabffabffab;
mem[3369] = 80'h0010ffabffabffabffab;
mem[3370] = 80'h0010ffabffabffabffab;
mem[3371] = 80'h0010ffabffabffabffab;
mem[3372] = 80'h0010ffabffabffabffab;
mem[3373] = 80'h0010ffabffabffabffab;
mem[3374] = 80'h0010ffabffabffabffab;
mem[3375] = 80'h0010ffabffabffabffab;
mem[3376] = 80'h0010ffabffabffabffab;
mem[3377] = 80'h0010ffabffabffabffab;
mem[3378] = 80'h0010ffabffabffabffab;
mem[3379] = 80'h0010ffabffabffabffab;
mem[3380] = 80'h0010ffabffabffabffab;
mem[3381] = 80'h0010ffabffabffabffab;
mem[3382] = 80'h0010ffabffabffabffab;
mem[3383] = 80'h0010ffabffabffabffab;
mem[3384] = 80'h0010ffabffabffabffab;
mem[3385] = 80'h0010ffabffabffabffab;
mem[3386] = 80'h0010ffabffabffabffab;
mem[3387] = 80'h0010ffabffabffabffab;
mem[3388] = 80'h0010ffabffabffabffab;
mem[3389] = 80'h0010ffabffabffabffab;
mem[3390] = 80'h0010ffabffabffabffab;
mem[3391] = 80'h0010ffabffabffabffab;
mem[3392] = 80'h0010ffabffabffabffab;
mem[3393] = 80'h0010ffabffabffabffab;
mem[3394] = 80'h0010ffabffabffabffab;
mem[3395] = 80'h0010ffabffabffabffab;
mem[3396] = 80'h0010ffabffabffabffab;
mem[3397] = 80'h0010ffabffabffabffab;
mem[3398] = 80'h0010ffabffabffabffab;
mem[3399] = 80'h0010ffabffabffabffab;
mem[3400] = 80'h0010ffabffabffabffab;
mem[3401] = 80'h0010ffabffabffabffab;
mem[3402] = 80'h0010ffabffabffabffab;
mem[3403] = 80'h0010ffabffabffabffab;
mem[3404] = 80'h0010ffabffabffabffab;
mem[3405] = 80'h0010ffabffabffabffab;
mem[3406] = 80'h0010ffabffabffabffab;
mem[3407] = 80'h0010ffabffabffabffab;
mem[3408] = 80'h0010ffabffabffabffab;
mem[3409] = 80'h0010ffabffabffabffab;
mem[3410] = 80'h0010ffabffabffabffab;
mem[3411] = 80'h0010ffabffabffabffab;
mem[3412] = 80'h0010ffabffabffabffab;
mem[3413] = 80'h0010ffabffabffabffab;
mem[3414] = 80'h0010ffabffabffabffab;
mem[3415] = 80'h0010ffabffabffabffab;
mem[3416] = 80'h0010ffabffabffabffab;
mem[3417] = 80'h0010ffabffabffabffab;
mem[3418] = 80'h0010ffabffabffabffab;
mem[3419] = 80'h0010ffabffabffabffab;
mem[3420] = 80'h0010ffabffabffabffab;
mem[3421] = 80'h0010ffabffabffabffab;
mem[3422] = 80'h0010ffabffabffabffab;
mem[3423] = 80'h0010ffabffabffabffab;
mem[3424] = 80'h0010ffabffabffabffab;
mem[3425] = 80'h0010ffabffabffabffab;
mem[3426] = 80'h0010ffabffabffabffab;
mem[3427] = 80'h0010ffabffabffabffab;
mem[3428] = 80'h0010ffabffabffabffab;
mem[3429] = 80'h0010ffabffabffabffab;
mem[3430] = 80'h0010ffabffabffabffab;
mem[3431] = 80'h0010ffabffabffabffab;
mem[3432] = 80'h0010ffabffabffabffab;
mem[3433] = 80'h0010ffabffabffabffab;
mem[3434] = 80'h0010ffabffabffabffab;
mem[3435] = 80'h0010ffabffabffabffab;
mem[3436] = 80'h0010ffabffabffabffab;
mem[3437] = 80'h0010ffabffabffabffab;
mem[3438] = 80'h0010ffabffabffabffab;
mem[3439] = 80'h0010ffabffabffabffab;
mem[3440] = 80'h0010ffabffabffabffab;
mem[3441] = 80'h0010ffabffabffabffab;
mem[3442] = 80'h0010ffabffabffabffab;
mem[3443] = 80'h0010ffabffabffabffab;
mem[3444] = 80'h0010ffabffabffabffab;
mem[3445] = 80'h0010ffabffabffabffab;
mem[3446] = 80'h0010ffabffabffabffab;
mem[3447] = 80'h0010ffabffabffabffab;
mem[3448] = 80'h0010ffabffabffabffab;
mem[3449] = 80'h0010ffabffabffabffab;
mem[3450] = 80'h0010ffabffabffabffab;
mem[3451] = 80'h0010ffabffabffabffab;
mem[3452] = 80'h0010ffabffabffabffab;
mem[3453] = 80'h0010ffabffabffabffab;
mem[3454] = 80'h0010ffabffabffabffab;
mem[3455] = 80'h0010ffabffabffabffab;
mem[3456] = 80'h0010ffabffabffabffab;
mem[3457] = 80'h0010ffabffabffabffab;
mem[3458] = 80'h0010ffabffabffabffab;
mem[3459] = 80'h0010ffabffabffabffab;
mem[3460] = 80'h0010ffabffabffabffab;
mem[3461] = 80'h0010ffabffabffabffab;
mem[3462] = 80'h0010ffabffabffabffab;
mem[3463] = 80'h0010ffabffabffabffab;
mem[3464] = 80'h0010ffabffabffabffab;
mem[3465] = 80'h0010ffabffabffabffab;
mem[3466] = 80'h0010ffabffabffabffab;
mem[3467] = 80'h0010ffabffabffabffab;
mem[3468] = 80'h0010ffabffabffabffab;
mem[3469] = 80'h0010ffabffabffabffab;
mem[3470] = 80'h0010ffabffabffabffab;
mem[3471] = 80'h0010ffabffabffabffab;
mem[3472] = 80'h0010ffabffabffabffab;
mem[3473] = 80'h0010ffabffabffabffab;
mem[3474] = 80'h0010ffabffabffabffab;
mem[3475] = 80'h0010ffabffabffabffab;
mem[3476] = 80'h0010ffabffabffabffab;
mem[3477] = 80'h0010ffabffabff44523f;
mem[3478] = 80'h001002e335d1c6840cc4;
mem[3479] = 80'h0010524936f083562cef;
mem[3480] = 80'h011568fcbbeeea000000;
mem[3481] = 80'h00000000000000000000;
mem[3482] = 80'h00000000000000000000;
mem[3483] = 80'h00000000000000000000;
mem[3484] = 80'h00000000000000000000;
mem[3485] = 80'h00000000000000000000;
mem[3486] = 80'h10100000010000010010;
mem[3487] = 80'h00109400000208004500;
mem[3488] = 80'h0010051489bc0000fffd;
mem[3489] = 80'h0010aad7c0550102c000;
mem[3490] = 80'h00100001ffabffabffab;
mem[3491] = 80'h0010ffabffabffabffab;
mem[3492] = 80'h0010ffabffabffabffab;
mem[3493] = 80'h0010ffabffabffabffab;
mem[3494] = 80'h0010ffabffabffabffab;
mem[3495] = 80'h0010ffabffabffabffab;
mem[3496] = 80'h0010ffabffabffabffab;
mem[3497] = 80'h0010ffabffabffabffab;
mem[3498] = 80'h0010ffabffabffabffab;
mem[3499] = 80'h0010ffabffabffabffab;
mem[3500] = 80'h0010ffabffabffabffab;
mem[3501] = 80'h0010ffabffabffabffab;
mem[3502] = 80'h0010ffabffabffabffab;
mem[3503] = 80'h0010ffabffabffabffab;
mem[3504] = 80'h0010ffabffabffabffab;
mem[3505] = 80'h0010ffabffabffabffab;
mem[3506] = 80'h0010ffabffabffabffab;
mem[3507] = 80'h0010ffabffabffabffab;
mem[3508] = 80'h0010ffabffabffabffab;
mem[3509] = 80'h0010ffabffabffabffab;
mem[3510] = 80'h0010ffabffabffabffab;
mem[3511] = 80'h0010ffabffabffabffab;
mem[3512] = 80'h0010ffabffabffabffab;
mem[3513] = 80'h0010ffabffabffabffab;
mem[3514] = 80'h0010ffabffabffabffab;
mem[3515] = 80'h0010ffabffabffabffab;
mem[3516] = 80'h0010ffabffabffabffab;
mem[3517] = 80'h0010ffabffabffabffab;
mem[3518] = 80'h0010ffabffabffabffab;
mem[3519] = 80'h0010ffabffabffabffab;
mem[3520] = 80'h0010ffabffabffabffab;
mem[3521] = 80'h0010ffabffabffabffab;
mem[3522] = 80'h0010ffabffabffabffab;
mem[3523] = 80'h0010ffabffabffabffab;
mem[3524] = 80'h0010ffabffabffabffab;
mem[3525] = 80'h0010ffabffabffabffab;
mem[3526] = 80'h0010ffabffabffabffab;
mem[3527] = 80'h0010ffabffabffabffab;
mem[3528] = 80'h0010ffabffabffabffab;
mem[3529] = 80'h0010ffabffabffabffab;
mem[3530] = 80'h0010ffabffabffabffab;
mem[3531] = 80'h0010ffabffabffabffab;
mem[3532] = 80'h0010ffabffabffabffab;
mem[3533] = 80'h0010ffabffabffabffab;
mem[3534] = 80'h0010ffabffabffabffab;
mem[3535] = 80'h0010ffabffabffabffab;
mem[3536] = 80'h0010ffabffabffabffab;
mem[3537] = 80'h0010ffabffabffabffab;
mem[3538] = 80'h0010ffabffabffabffab;
mem[3539] = 80'h0010ffabffabffabffab;
mem[3540] = 80'h0010ffabffabffabffab;
mem[3541] = 80'h0010ffabffabffabffab;
mem[3542] = 80'h0010ffabffabffabffab;
mem[3543] = 80'h0010ffabffabffabffab;
mem[3544] = 80'h0010ffabffabffabffab;
mem[3545] = 80'h0010ffabffabffabffab;
mem[3546] = 80'h0010ffabffabffabffab;
mem[3547] = 80'h0010ffabffabffabffab;
mem[3548] = 80'h0010ffabffabffabffab;
mem[3549] = 80'h0010ffabffabffabffab;
mem[3550] = 80'h0010ffabffabffabffab;
mem[3551] = 80'h0010ffabffabffabffab;
mem[3552] = 80'h0010ffabffabffabffab;
mem[3553] = 80'h0010ffabffabffabffab;
mem[3554] = 80'h0010ffabffabffabffab;
mem[3555] = 80'h0010ffabffabffabffab;
mem[3556] = 80'h0010ffabffabffabffab;
mem[3557] = 80'h0010ffabffabffabffab;
mem[3558] = 80'h0010ffabffabffabffab;
mem[3559] = 80'h0010ffabffabffabffab;
mem[3560] = 80'h0010ffabffabffabffab;
mem[3561] = 80'h0010ffabffabffabffab;
mem[3562] = 80'h0010ffabffabffabffab;
mem[3563] = 80'h0010ffabffabffabffab;
mem[3564] = 80'h0010ffabffabffabffab;
mem[3565] = 80'h0010ffabffabffabffab;
mem[3566] = 80'h0010ffabffabffabffab;
mem[3567] = 80'h0010ffabffabffabffab;
mem[3568] = 80'h0010ffabffabffabffab;
mem[3569] = 80'h0010ffabffabffabffab;
mem[3570] = 80'h0010ffabffabffabffab;
mem[3571] = 80'h0010ffabffabffabffab;
mem[3572] = 80'h0010ffabffabffabffab;
mem[3573] = 80'h0010ffabffabffabffab;
mem[3574] = 80'h0010ffabffabffabffab;
mem[3575] = 80'h0010ffabffabffabffab;
mem[3576] = 80'h0010ffabffabffabffab;
mem[3577] = 80'h0010ffabffabffabffab;
mem[3578] = 80'h0010ffabffabffabffab;
mem[3579] = 80'h0010ffabffabffabffab;
mem[3580] = 80'h0010ffabffabffabffab;
mem[3581] = 80'h0010ffabffabffabffab;
mem[3582] = 80'h0010ffabffabffabffab;
mem[3583] = 80'h0010ffabffabffabffab;
mem[3584] = 80'h0010ffabffabffabffab;
mem[3585] = 80'h0010ffabffabffabffab;
mem[3586] = 80'h0010ffabffabffabffab;
mem[3587] = 80'h0010ffabffabffabffab;
mem[3588] = 80'h0010ffabffabffabffab;
mem[3589] = 80'h0010ffabffabffabffab;
mem[3590] = 80'h0010ffabffabffabffab;
mem[3591] = 80'h0010ffabffabffabffab;
mem[3592] = 80'h0010ffabffabffabffab;
mem[3593] = 80'h0010ffabffabffabffab;
mem[3594] = 80'h0010ffabffabffabffab;
mem[3595] = 80'h0010ffabffabffabffab;
mem[3596] = 80'h0010ffabffabffabffab;
mem[3597] = 80'h0010ffabffabffabffab;
mem[3598] = 80'h0010ffabffabffabffab;
mem[3599] = 80'h0010ffabffabffabffab;
mem[3600] = 80'h0010ffabffabffabffab;
mem[3601] = 80'h0010ffabffabffabffab;
mem[3602] = 80'h0010ffabffabffabffab;
mem[3603] = 80'h0010ffabffabffabffab;
mem[3604] = 80'h0010ffabffabffabffab;
mem[3605] = 80'h0010ffabffabffabffab;
mem[3606] = 80'h0010ffabffabffabffab;
mem[3607] = 80'h0010ffabffabffabffab;
mem[3608] = 80'h0010ffabffabffabffab;
mem[3609] = 80'h0010ffabffabffabffab;
mem[3610] = 80'h0010ffabffabffabffab;
mem[3611] = 80'h0010ffabffabffabffab;
mem[3612] = 80'h0010ffabffabffabffab;
mem[3613] = 80'h0010ffabffabffabffab;
mem[3614] = 80'h0010ffabffabffabffab;
mem[3615] = 80'h0010ffabffabffabffab;
mem[3616] = 80'h0010ffabffabffabffab;
mem[3617] = 80'h0010ffabffabffabffab;
mem[3618] = 80'h0010ffabffabffabffab;
mem[3619] = 80'h0010ffabffabffabffab;
mem[3620] = 80'h0010ffabffabffabffab;
mem[3621] = 80'h0010ffabffabffabffab;
mem[3622] = 80'h0010ffabffabffabffab;
mem[3623] = 80'h0010ffabffabffabffab;
mem[3624] = 80'h0010ffabffabffabffab;
mem[3625] = 80'h0010ffabffabffabffab;
mem[3626] = 80'h0010ffabffabffabffab;
mem[3627] = 80'h0010ffabffabffabffab;
mem[3628] = 80'h0010ffabffabffabffab;
mem[3629] = 80'h0010ffabffabffabffab;
mem[3630] = 80'h0010ffabffabffabffab;
mem[3631] = 80'h0010ffabffabffabffab;
mem[3632] = 80'h0010ffabffabffabffab;
mem[3633] = 80'h0010ffabffabffabffab;
mem[3634] = 80'h0010ffabffabffabffab;
mem[3635] = 80'h0010ffabffabffabffab;
mem[3636] = 80'h0010ffabffabffabffab;
mem[3637] = 80'h0010ffabffabffabffab;
mem[3638] = 80'h0010ffabffabffabffab;
mem[3639] = 80'h0010ffabffabffabffab;
mem[3640] = 80'h0010ffabffabffabffab;
mem[3641] = 80'h0010ffabffabffabffab;
mem[3642] = 80'h0010ffabffabffabffab;
mem[3643] = 80'h0010ffabffabffabffab;
mem[3644] = 80'h0010ffabffabffabffab;
mem[3645] = 80'h0010ffabffabffabffab;
mem[3646] = 80'h0010ffabffabffabffab;
mem[3647] = 80'h0010ffabffabffab4376;
mem[3648] = 80'h0010fbe832215e463ce3;
mem[3649] = 80'h0010d53e75d01366d302;
mem[3650] = 80'h0116c1dd0cd6b9300000;
mem[3651] = 80'h10100000010000010010;
mem[3652] = 80'h00109400000208004500;
mem[3653] = 80'h0010029f89bd0000fffd;
mem[3654] = 80'h0010ad4bc0550102c000;
mem[3655] = 80'h00100001ffabffabffab;
mem[3656] = 80'h0010ffabffabffabffab;
mem[3657] = 80'h0010ffabffabffabffab;
mem[3658] = 80'h0010ffabffabffabffab;
mem[3659] = 80'h0010ffabffabffabffab;
mem[3660] = 80'h0010ffabffabffabffab;
mem[3661] = 80'h0010ffabffabffabffab;
mem[3662] = 80'h0010ffabffabffabffab;
mem[3663] = 80'h0010ffabffabffabffab;
mem[3664] = 80'h0010ffabffabffabffab;
mem[3665] = 80'h0010ffabffabffabffab;
mem[3666] = 80'h0010ffabffabffabffab;
mem[3667] = 80'h0010ffabffabffabffab;
mem[3668] = 80'h0010ffabffabffabffab;
mem[3669] = 80'h0010ffabffabffabffab;
mem[3670] = 80'h0010ffabffabffabffab;
mem[3671] = 80'h0010ffabffabffabffab;
mem[3672] = 80'h0010ffabffabffabffab;
mem[3673] = 80'h0010ffabffabffabffab;
mem[3674] = 80'h0010ffabffabffabffab;
mem[3675] = 80'h0010ffabffabffabffab;
mem[3676] = 80'h0010ffabffabffabffab;
mem[3677] = 80'h0010ffabffabffabffab;
mem[3678] = 80'h0010ffabffabffabffab;
mem[3679] = 80'h0010ffabffabffabffab;
mem[3680] = 80'h0010ffabffabffabffab;
mem[3681] = 80'h0010ffabffabffabffab;
mem[3682] = 80'h0010ffabffabffabffab;
mem[3683] = 80'h0010ffabffabffabffab;
mem[3684] = 80'h0010ffabffabffabffab;
mem[3685] = 80'h0010ffabffabffabffab;
mem[3686] = 80'h0010ffabffabffabffab;
mem[3687] = 80'h0010ffabffabffabffab;
mem[3688] = 80'h0010ffabffabffabffab;
mem[3689] = 80'h0010ffabffabffabffab;
mem[3690] = 80'h0010ffabffabffabffab;
mem[3691] = 80'h0010ffabffabffabffab;
mem[3692] = 80'h0010ffabffabffabffab;
mem[3693] = 80'h0010ffabffabffabffab;
mem[3694] = 80'h0010ffabffabffabffab;
mem[3695] = 80'h0010ffabffabffabffab;
mem[3696] = 80'h0010ffabffabffabffab;
mem[3697] = 80'h0010ffabffabffabffab;
mem[3698] = 80'h0010ffabffabffabffab;
mem[3699] = 80'h0010ffabffabffabffab;
mem[3700] = 80'h0010ffabffabffabffab;
mem[3701] = 80'h0010ffabffabffabffab;
mem[3702] = 80'h0010ffabffabffabffab;
mem[3703] = 80'h0010ffabffabffabffab;
mem[3704] = 80'h0010ffabffabffabffab;
mem[3705] = 80'h0010ffabffabffabffab;
mem[3706] = 80'h0010ffabffabffabffab;
mem[3707] = 80'h0010ffabffabffabffab;
mem[3708] = 80'h0010ffabffabffabffab;
mem[3709] = 80'h0010ffabffabffabffab;
mem[3710] = 80'h0010ffabffabffabffab;
mem[3711] = 80'h0010ffabffabffabffab;
mem[3712] = 80'h0010ffabffabffabffab;
mem[3713] = 80'h0010ffabffabffabffab;
mem[3714] = 80'h0010ffabffabffabffab;
mem[3715] = 80'h0010ffabffabffabffab;
mem[3716] = 80'h0010ffabffabffabffab;
mem[3717] = 80'h0010ffabffabffabffab;
mem[3718] = 80'h0010ffabffabffabffab;
mem[3719] = 80'h0010ffabffabffabffab;
mem[3720] = 80'h0010ffabffabffabffab;
mem[3721] = 80'h0010ffabffabffabffab;
mem[3722] = 80'h0010ffabffabffabffab;
mem[3723] = 80'h0010ffabffabffabffab;
mem[3724] = 80'h0010ffabffabffabffab;
mem[3725] = 80'h0010ffabffabffabffab;
mem[3726] = 80'h0010ffabffabffabffab;
mem[3727] = 80'h0010ffabffabffabffab;
mem[3728] = 80'h0010ffabffabffabffab;
mem[3729] = 80'h0010ffabffabffabffab;
mem[3730] = 80'h0010ffabffabffabffab;
mem[3731] = 80'h0010ffabffabffabffab;
mem[3732] = 80'h0010ffabffabffabffab;
mem[3733] = 80'h0010ffabffabffabffab;
mem[3734] = 80'h0010ff420725c4ea589c;
mem[3735] = 80'h0010f9f73152d38002a5;
mem[3736] = 80'h0010377803299f729642;
mem[3737] = 80'h01112200000000000000;
mem[3738] = 80'h10100000010000010010;
mem[3739] = 80'h00109400000208004500;
mem[3740] = 80'h0010016689be0000fffd;
mem[3741] = 80'h0010ae83c0550102c000;
mem[3742] = 80'h00100001ffabffabffab;
mem[3743] = 80'h0010ffabffabffabffab;
mem[3744] = 80'h0010ffabffabffabffab;
mem[3745] = 80'h0010ffabffabffabffab;
mem[3746] = 80'h0010ffabffabffabffab;
mem[3747] = 80'h0010ffabffabffabffab;
mem[3748] = 80'h0010ffabffabffabffab;
mem[3749] = 80'h0010ffabffabffabffab;
mem[3750] = 80'h0010ffabffabffabffab;
mem[3751] = 80'h0010ffabffabffabffab;
mem[3752] = 80'h0010ffabffabffabffab;
mem[3753] = 80'h0010ffabffabffabffab;
mem[3754] = 80'h0010ffabffabffabffab;
mem[3755] = 80'h0010ffabffabffabffab;
mem[3756] = 80'h0010ffabffabffabffab;
mem[3757] = 80'h0010ffabffabffabffab;
mem[3758] = 80'h0010ffabffabffabffab;
mem[3759] = 80'h0010ffabffabffabffab;
mem[3760] = 80'h0010ffabffabffabffab;
mem[3761] = 80'h0010ffabffabffabffab;
mem[3762] = 80'h0010ffabffabffabffab;
mem[3763] = 80'h0010ffabffabffabffab;
mem[3764] = 80'h0010ffabffabffabffab;
mem[3765] = 80'h0010ffabffabffabffab;
mem[3766] = 80'h0010ffabffabffabffab;
mem[3767] = 80'h0010ffabffabffabffab;
mem[3768] = 80'h0010ffabffabffabffab;
mem[3769] = 80'h0010ffabffabffabffab;
mem[3770] = 80'h0010ffabffabffabffab;
mem[3771] = 80'h0010ffabffabffabffab;
mem[3772] = 80'h0010ffabffabffabffab;
mem[3773] = 80'h0010ffabffabffabffab;
mem[3774] = 80'h0010ffabffabffabffab;
mem[3775] = 80'h0010ffabffabffabffab;
mem[3776] = 80'h0010ffabffabffabffab;
mem[3777] = 80'h0010ffabffabffabffab;
mem[3778] = 80'h0010ffabffabffabffab;
mem[3779] = 80'h0010ffabffabffabffab;
mem[3780] = 80'h0010ffabffabffabffab;
mem[3781] = 80'h0010ffabffabffabffab;
mem[3782] = 80'h0010419547b182d2db39;
mem[3783] = 80'h0010ab46dae59e7366c5;
mem[3784] = 80'h01108e4bfefb382d9898;
mem[3785] = 80'h10100000010000010010;
mem[3786] = 80'h00109400000208004500;
mem[3787] = 80'h001003a389bf0000fffd;
mem[3788] = 80'h0010ac45c0550102c000;
mem[3789] = 80'h00100001ffabffabffab;
mem[3790] = 80'h0010ffabffabffabffab;
mem[3791] = 80'h0010ffabffabffabffab;
mem[3792] = 80'h0010ffabffabffabffab;
mem[3793] = 80'h0010ffabffabffabffab;
mem[3794] = 80'h0010ffabffabffabffab;
mem[3795] = 80'h0010ffabffabffabffab;
mem[3796] = 80'h0010ffabffabffabffab;
mem[3797] = 80'h0010ffabffabffabffab;
mem[3798] = 80'h0010ffabffabffabffab;
mem[3799] = 80'h0010ffabffabffabffab;
mem[3800] = 80'h0010ffabffabffabffab;
mem[3801] = 80'h0010ffabffabffabffab;
mem[3802] = 80'h0010ffabffabffabffab;
mem[3803] = 80'h0010ffabffabffabffab;
mem[3804] = 80'h0010ffabffabffabffab;
mem[3805] = 80'h0010ffabffabffabffab;
mem[3806] = 80'h0010ffabffabffabffab;
mem[3807] = 80'h0010ffabffabffabffab;
mem[3808] = 80'h0010ffabffabffabffab;
mem[3809] = 80'h0010ffabffabffabffab;
mem[3810] = 80'h0010ffabffabffabffab;
mem[3811] = 80'h0010ffabffabffabffab;
mem[3812] = 80'h0010ffabffabffabffab;
mem[3813] = 80'h0010ffabffabffabffab;
mem[3814] = 80'h0010ffabffabffabffab;
mem[3815] = 80'h0010ffabffabffabffab;
mem[3816] = 80'h0010ffabffabffabffab;
mem[3817] = 80'h0010ffabffabffabffab;
mem[3818] = 80'h0010ffabffabffabffab;
mem[3819] = 80'h0010ffabffabffabffab;
mem[3820] = 80'h0010ffabffabffabffab;
mem[3821] = 80'h0010ffabffabffabffab;
mem[3822] = 80'h0010ffabffabffabffab;
mem[3823] = 80'h0010ffabffabffabffab;
mem[3824] = 80'h0010ffabffabffabffab;
mem[3825] = 80'h0010ffabffabffabffab;
mem[3826] = 80'h0010ffabffabffabffab;
mem[3827] = 80'h0010ffabffabffabffab;
mem[3828] = 80'h0010ffabffabffabffab;
mem[3829] = 80'h0010ffabffabffabffab;
mem[3830] = 80'h0010ffabffabffabffab;
mem[3831] = 80'h0010ffabffabffabffab;
mem[3832] = 80'h0010ffabffabffabffab;
mem[3833] = 80'h0010ffabffabffabffab;
mem[3834] = 80'h0010ffabffabffabffab;
mem[3835] = 80'h0010ffabffabffabffab;
mem[3836] = 80'h0010ffabffabffabffab;
mem[3837] = 80'h0010ffabffabffabffab;
mem[3838] = 80'h0010ffabffabffabffab;
mem[3839] = 80'h0010ffabffabffabffab;
mem[3840] = 80'h0010ffabffabffabffab;
mem[3841] = 80'h0010ffabffabffabffab;
mem[3842] = 80'h0010ffabffabffabffab;
mem[3843] = 80'h0010ffabffabffabffab;
mem[3844] = 80'h0010ffabffabffabffab;
mem[3845] = 80'h0010ffabffabffabffab;
mem[3846] = 80'h0010ffabffabffabffab;
mem[3847] = 80'h0010ffabffabffabffab;
mem[3848] = 80'h0010ffabffabffabffab;
mem[3849] = 80'h0010ffabffabffabffab;
mem[3850] = 80'h0010ffabffabffabffab;
mem[3851] = 80'h0010ffabffabffabffab;
mem[3852] = 80'h0010ffabffabffabffab;
mem[3853] = 80'h0010ffabffabffabffab;
mem[3854] = 80'h0010ffabffabffabffab;
mem[3855] = 80'h0010ffabffabffabffab;
mem[3856] = 80'h0010ffabffabffabffab;
mem[3857] = 80'h0010ffabffabffabffab;
mem[3858] = 80'h0010ffabffabffabffab;
mem[3859] = 80'h0010ffabffabffabffab;
mem[3860] = 80'h0010ffabffabffabffab;
mem[3861] = 80'h0010ffabffabffabffab;
mem[3862] = 80'h0010ffabffabffabffab;
mem[3863] = 80'h0010ffabffabffabffab;
mem[3864] = 80'h0010ffabffabffabffab;
mem[3865] = 80'h0010ffabffabffabffab;
mem[3866] = 80'h0010ffabffabffabffab;
mem[3867] = 80'h0010ffabffabffabffab;
mem[3868] = 80'h0010ffabffabffabffab;
mem[3869] = 80'h0010ffabffabffabffab;
mem[3870] = 80'h0010ffabffabffabffab;
mem[3871] = 80'h0010ffabffabffabffab;
mem[3872] = 80'h0010ffabffabffabffab;
mem[3873] = 80'h0010ffabffabffabffab;
mem[3874] = 80'h0010ffabffabffabffab;
mem[3875] = 80'h0010ffabffabffabffab;
mem[3876] = 80'h0010ffabffabffabffab;
mem[3877] = 80'h0010ffabffabffabffab;
mem[3878] = 80'h0010ffabffabffabffab;
mem[3879] = 80'h0010ffabffabffabffab;
mem[3880] = 80'h0010ffabffabffabffab;
mem[3881] = 80'h0010ffabffabffabffab;
mem[3882] = 80'h0010ffabffabffabffab;
mem[3883] = 80'h0010ffabffabffabffab;
mem[3884] = 80'h0010ffabffabffabffab;
mem[3885] = 80'h0010ffabffabffabffab;
mem[3886] = 80'h0010ffabffabffabffab;
mem[3887] = 80'h0010ffabffabffabffab;
mem[3888] = 80'h0010ffabffabffabffab;
mem[3889] = 80'h0010ffabffabffabffab;
mem[3890] = 80'h0010ffabffabffabffab;
mem[3891] = 80'h0010ffabffabffabffab;
mem[3892] = 80'h0010ffabffabffabffab;
mem[3893] = 80'h0010ffabffabffabffab;
mem[3894] = 80'h0010ffabffabffabffab;
mem[3895] = 80'h0010ffabffabffabffab;
mem[3896] = 80'h0010ffabffabffabffab;
mem[3897] = 80'h0010ffabffabffabffab;
mem[3898] = 80'h0010ffabffabffabffab;
mem[3899] = 80'h0010ffabffabffabffab;
mem[3900] = 80'h0010ffabffabff40e499;
mem[3901] = 80'h00109d5aab198660945d;
mem[3902] = 80'h0010086ba3839410c6f3;
mem[3903] = 80'h0115b109e0d2dc000000;
mem[3904] = 80'h10100000010000010010;
mem[3905] = 80'h00109400000208004500;
mem[3906] = 80'h001004be89c00000fffd;
mem[3907] = 80'h0010ab29c0550102c000;
mem[3908] = 80'h00100001ffabffabffab;
mem[3909] = 80'h0010ffabffabffabffab;
mem[3910] = 80'h0010ffabffabffabffab;
mem[3911] = 80'h0010ffabffabffabffab;
mem[3912] = 80'h0010ffabffabffabffab;
mem[3913] = 80'h0010ffabffabffabffab;
mem[3914] = 80'h0010ffabffabffabffab;
mem[3915] = 80'h0010ffabffabffabffab;
mem[3916] = 80'h0010ffabffabffabffab;
mem[3917] = 80'h0010ffabffabffabffab;
mem[3918] = 80'h0010ffabffabffabffab;
mem[3919] = 80'h0010ffabffabffabffab;
mem[3920] = 80'h0010ffabffabffabffab;
mem[3921] = 80'h0010ffabffabffabffab;
mem[3922] = 80'h0010ffabffabffabffab;
mem[3923] = 80'h0010ffabffabffabffab;
mem[3924] = 80'h0010ffabffabffabffab;
mem[3925] = 80'h0010ffabffabffabffab;
mem[3926] = 80'h0010ffabffabffabffab;
mem[3927] = 80'h0010ffabffabffabffab;
mem[3928] = 80'h0010ffabffabffabffab;
mem[3929] = 80'h0010ffabffabffabffab;
mem[3930] = 80'h0010ffabffabffabffab;
mem[3931] = 80'h0010ffabffabffabffab;
mem[3932] = 80'h0010ffabffabffabffab;
mem[3933] = 80'h0010ffabffabffabffab;
mem[3934] = 80'h0010ffabffabffabffab;
mem[3935] = 80'h0010ffabffabffabffab;
mem[3936] = 80'h0010ffabffabffabffab;
mem[3937] = 80'h0010ffabffabffabffab;
mem[3938] = 80'h0010ffabffabffabffab;
mem[3939] = 80'h0010ffabffabffabffab;
mem[3940] = 80'h0010ffabffabffabffab;
mem[3941] = 80'h0010ffabffabffabffab;
mem[3942] = 80'h0010ffabffabffabffab;
mem[3943] = 80'h0010ffabffabffabffab;
mem[3944] = 80'h0010ffabffabffabffab;
mem[3945] = 80'h0010ffabffabffabffab;
mem[3946] = 80'h0010ffabffabffabffab;
mem[3947] = 80'h0010ffabffabffabffab;
mem[3948] = 80'h0010ffabffabffabffab;
mem[3949] = 80'h0010ffabffabffabffab;
mem[3950] = 80'h0010ffabffabffabffab;
mem[3951] = 80'h0010ffabffabffabffab;
mem[3952] = 80'h0010ffabffabffabffab;
mem[3953] = 80'h0010ffabffabffabffab;
mem[3954] = 80'h0010ffabffabffabffab;
mem[3955] = 80'h0010ffabffabffabffab;
mem[3956] = 80'h0010ffabffabffabffab;
mem[3957] = 80'h0010ffabffabffabffab;
mem[3958] = 80'h0010ffabffabffabffab;
mem[3959] = 80'h0010ffabffabffabffab;
mem[3960] = 80'h0010ffabffabffabffab;
mem[3961] = 80'h0010ffabffabffabffab;
mem[3962] = 80'h0010ffabffabffabffab;
mem[3963] = 80'h0010ffabffabffabffab;
mem[3964] = 80'h0010ffabffabffabffab;
mem[3965] = 80'h0010ffabffabffabffab;
mem[3966] = 80'h0010ffabffabffabffab;
mem[3967] = 80'h0010ffabffabffabffab;
mem[3968] = 80'h0010ffabffabffabffab;
mem[3969] = 80'h0010ffabffabffabffab;
mem[3970] = 80'h0010ffabffabffabffab;
mem[3971] = 80'h0010ffabffabffabffab;
mem[3972] = 80'h0010ffabffabffabffab;
mem[3973] = 80'h0010ffabffabffabffab;
mem[3974] = 80'h0010ffabffabffabffab;
mem[3975] = 80'h0010ffabffabffabffab;
mem[3976] = 80'h0010ffabffabffabffab;
mem[3977] = 80'h0010ffabffabffabffab;
mem[3978] = 80'h0010ffabffabffabffab;
mem[3979] = 80'h0010ffabffabffabffab;
mem[3980] = 80'h0010ffabffabffabffab;
mem[3981] = 80'h0010ffabffabffabffab;
mem[3982] = 80'h0010ffabffabffabffab;
mem[3983] = 80'h0010ffabffabffabffab;
mem[3984] = 80'h0010ffabffabffabffab;
mem[3985] = 80'h0010ffabffabffabffab;
mem[3986] = 80'h0010ffabffabffabffab;
mem[3987] = 80'h0010ffabffabffabffab;
mem[3988] = 80'h0010ffabffabffabffab;
mem[3989] = 80'h0010ffabffabffabffab;
mem[3990] = 80'h0010ffabffabffabffab;
mem[3991] = 80'h0010ffabffabffabffab;
mem[3992] = 80'h0010ffabffabffabffab;
mem[3993] = 80'h0010ffabffabffabffab;
mem[3994] = 80'h0010ffabffabffabffab;
mem[3995] = 80'h0010ffabffabffabffab;
mem[3996] = 80'h0010ffabffabffabffab;
mem[3997] = 80'h0010ffabffabffabffab;
mem[3998] = 80'h0010ffabffabffabffab;
mem[3999] = 80'h0010ffabffabffabffab;
mem[4000] = 80'h0010ffabffabffabffab;
mem[4001] = 80'h0010ffabffabffabffab;
mem[4002] = 80'h0010ffabffabffabffab;
mem[4003] = 80'h0010ffabffabffabffab;
mem[4004] = 80'h0010ffabffabffabffab;
mem[4005] = 80'h0010ffabffabffabffab;
mem[4006] = 80'h0010ffabffabffabffab;
mem[4007] = 80'h0010ffabffabffabffab;
mem[4008] = 80'h0010ffabffabffabffab;
mem[4009] = 80'h0010ffabffabffabffab;
mem[4010] = 80'h0010ffabffabffabffab;
mem[4011] = 80'h0010ffabffabffabffab;
mem[4012] = 80'h0010ffabffabffabffab;
mem[4013] = 80'h0010ffabffabffabffab;
mem[4014] = 80'h0010ffabffabffabffab;
mem[4015] = 80'h0010ffabffabffabffab;
mem[4016] = 80'h0010ffabffabffabffab;
mem[4017] = 80'h0010ffabffabffabffab;
mem[4018] = 80'h0010ffabffabffabffab;
mem[4019] = 80'h0010ffabffabffabffab;
mem[4020] = 80'h0010ffabffabffabffab;
mem[4021] = 80'h0010ffabffabffabffab;
mem[4022] = 80'h0010ffabffabffabffab;
mem[4023] = 80'h0010ffabffabffabffab;
mem[4024] = 80'h0010ffabffabffabffab;
mem[4025] = 80'h0010ffabffabffabffab;
mem[4026] = 80'h0010ffabffabffabffab;
mem[4027] = 80'h0010ffabffabffabffab;
mem[4028] = 80'h0010ffabffabffabffab;
mem[4029] = 80'h0010ffabffabffabffab;
mem[4030] = 80'h0010ffabffabffabffab;
mem[4031] = 80'h0010ffabffabffabffab;
mem[4032] = 80'h0010ffabffabffabffab;
mem[4033] = 80'h0010ffabffabffabffab;
mem[4034] = 80'h0010ffabffabffabffab;
mem[4035] = 80'h0010ffabffabffabffab;
mem[4036] = 80'h0010ffabffabffabffab;
mem[4037] = 80'h0010ffabffabffabffab;
mem[4038] = 80'h0010ffabffabffabffab;
mem[4039] = 80'h0010ffabffabffabffab;
mem[4040] = 80'h0010ffabffabffabffab;
mem[4041] = 80'h0010ffabffabffabffab;
mem[4042] = 80'h0010ffabffabffabffab;
mem[4043] = 80'h0010ffabffabffabffab;
mem[4044] = 80'h0010ffabffabffabffab;
mem[4045] = 80'h0010ffabffabffabffab;
mem[4046] = 80'h0010ffabffabffabffab;
mem[4047] = 80'h0010ffabffabffabffab;
mem[4048] = 80'h0010ffabffabffabffab;
mem[4049] = 80'h0010ffabffabffabffab;
mem[4050] = 80'h0010ffabffabffabffab;
mem[4051] = 80'h0010ffabffabffabffab;
mem[4052] = 80'h0010ffabffabffabffab;
mem[4053] = 80'h0010ffabffabffabffab;
mem[4054] = 80'h0010ffabffabffabffab;
mem[4055] = 80'h00103f733c908140b94c;
mem[4056] = 80'h0010c3cce325c27b1bf3;
mem[4057] = 80'h0110e969daa3d6ce3e2e;
mem[4058] = 80'h00000000000000000000;
mem[4059] = 80'h00000000000000000000;
mem[4060] = 80'h00000000000000000000;
mem[4061] = 80'h00000000000000000000;
mem[4062] = 80'h00000000000000000000;
mem[4063] = 80'h00000000000000000000;
mem[4064] = 80'h00000000000000000000;
mem[4065] = 80'h00000000000000000000;
mem[4066] = 80'h00000000000000000000;
mem[4067] = 80'h00000000000000000000;
mem[4068] = 80'h00000000000000000000;
mem[4069] = 80'h00000000000000000000;
mem[4070] = 80'h00000000000000000000;
mem[4071] = 80'h00000000000000000000;
mem[4072] = 80'h00000000000000000000;
mem[4073] = 80'h00000000000000000000;
mem[4074] = 80'h00000000000000000000;
mem[4075] = 80'h00000000000000000000;
mem[4076] = 80'h00000000000000000000;
mem[4077] = 80'h10100000010000010010;
mem[4078] = 80'h00109400000208004500;
mem[4079] = 80'h0010054d89c10000fffd;
mem[4080] = 80'h0010aa99c0550102c000;
mem[4081] = 80'h00100001ffabffabffab;
mem[4082] = 80'h0010ffabffabffabffab;
mem[4083] = 80'h0010ffabffabffabffab;
mem[4084] = 80'h0010ffabffabffabffab;
mem[4085] = 80'h0010ffabffabffabffab;
mem[4086] = 80'h0010ffabffabffabffab;
mem[4087] = 80'h0010ffabffabffabffab;
mem[4088] = 80'h0010ffabffabffabffab;
mem[4089] = 80'h0010ffabffabffabffab;
mem[4090] = 80'h0010ffabffabffabffab;
mem[4091] = 80'h0010ffabffabffabffab;
mem[4092] = 80'h0010ffabffabffabffab;
mem[4093] = 80'h0010ffabffabffabffab;
mem[4094] = 80'h0010ffabffabffabffab;
mem[4095] = 80'h0010ffabffabffabffab;
mem[4096] = 80'h0010ffabffabffabffab;
mem[4097] = 80'h0010ffabffabffabffab;
mem[4098] = 80'h0010ffabffabffabffab;
mem[4099] = 80'h0010ffabffabffabffab;
mem[4100] = 80'h0010ffabffabffabffab;
mem[4101] = 80'h0010ffabffabffabffab;
mem[4102] = 80'h0010ffabffabffabffab;
mem[4103] = 80'h0010ffabffabffabffab;
mem[4104] = 80'h0010ffabffabffabffab;
mem[4105] = 80'h0010ffabffabffabffab;
mem[4106] = 80'h0010ffabffabffabffab;
mem[4107] = 80'h0010ffabffabffabffab;
mem[4108] = 80'h0010ffabffabffabffab;
mem[4109] = 80'h0010ffabffabffabffab;
mem[4110] = 80'h0010ffabffabffabffab;
mem[4111] = 80'h0010ffabffabffabffab;
mem[4112] = 80'h0010ffabffabffabffab;
mem[4113] = 80'h0010ffabffabffabffab;
mem[4114] = 80'h0010ffabffabffabffab;
mem[4115] = 80'h0010ffabffabffabffab;
mem[4116] = 80'h0010ffabffabffabffab;
mem[4117] = 80'h0010ffabffabffabffab;
mem[4118] = 80'h0010ffabffabffabffab;
mem[4119] = 80'h0010ffabffabffabffab;
mem[4120] = 80'h0010ffabffabffabffab;
mem[4121] = 80'h0010ffabffabffabffab;
mem[4122] = 80'h0010ffabffabffabffab;
mem[4123] = 80'h0010ffabffabffabffab;
mem[4124] = 80'h0010ffabffabffabffab;
mem[4125] = 80'h0010ffabffabffabffab;
mem[4126] = 80'h0010ffabffabffabffab;
mem[4127] = 80'h0010ffabffabffabffab;
mem[4128] = 80'h0010ffabffabffabffab;
mem[4129] = 80'h0010ffabffabffabffab;
mem[4130] = 80'h0010ffabffabffabffab;
mem[4131] = 80'h0010ffabffabffabffab;
mem[4132] = 80'h0010ffabffabffabffab;
mem[4133] = 80'h0010ffabffabffabffab;
mem[4134] = 80'h0010ffabffabffabffab;
mem[4135] = 80'h0010ffabffabffabffab;
mem[4136] = 80'h0010ffabffabffabffab;
mem[4137] = 80'h0010ffabffabffabffab;
mem[4138] = 80'h0010ffabffabffabffab;
mem[4139] = 80'h0010ffabffabffabffab;
mem[4140] = 80'h0010ffabffabffabffab;
mem[4141] = 80'h0010ffabffabffabffab;
mem[4142] = 80'h0010ffabffabffabffab;
mem[4143] = 80'h0010ffabffabffabffab;
mem[4144] = 80'h0010ffabffabffabffab;
mem[4145] = 80'h0010ffabffabffabffab;
mem[4146] = 80'h0010ffabffabffabffab;
mem[4147] = 80'h0010ffabffabffabffab;
mem[4148] = 80'h0010ffabffabffabffab;
mem[4149] = 80'h0010ffabffabffabffab;
mem[4150] = 80'h0010ffabffabffabffab;
mem[4151] = 80'h0010ffabffabffabffab;
mem[4152] = 80'h0010ffabffabffabffab;
mem[4153] = 80'h0010ffabffabffabffab;
mem[4154] = 80'h0010ffabffabffabffab;
mem[4155] = 80'h0010ffabffabffabffab;
mem[4156] = 80'h0010ffabffabffabffab;
mem[4157] = 80'h0010ffabffabffabffab;
mem[4158] = 80'h0010ffabffabffabffab;
mem[4159] = 80'h0010ffabffabffabffab;
mem[4160] = 80'h0010ffabffabffabffab;
mem[4161] = 80'h0010ffabffabffabffab;
mem[4162] = 80'h0010ffabffabffabffab;
mem[4163] = 80'h0010ffabffabffabffab;
mem[4164] = 80'h0010ffabffabffabffab;
mem[4165] = 80'h0010ffabffabffabffab;
mem[4166] = 80'h0010ffabffabffabffab;
mem[4167] = 80'h0010ffabffabffabffab;
mem[4168] = 80'h0010ffabffabffabffab;
mem[4169] = 80'h0010ffabffabffabffab;
mem[4170] = 80'h0010ffabffabffabffab;
mem[4171] = 80'h0010ffabffabffabffab;
mem[4172] = 80'h0010ffabffabffabffab;
mem[4173] = 80'h0010ffabffabffabffab;
mem[4174] = 80'h0010ffabffabffabffab;
mem[4175] = 80'h0010ffabffabffabffab;
mem[4176] = 80'h0010ffabffabffabffab;
mem[4177] = 80'h0010ffabffabffabffab;
mem[4178] = 80'h0010ffabffabffabffab;
mem[4179] = 80'h0010ffabffabffabffab;
mem[4180] = 80'h0010ffabffabffabffab;
mem[4181] = 80'h0010ffabffabffabffab;
mem[4182] = 80'h0010ffabffabffabffab;
mem[4183] = 80'h0010ffabffabffabffab;
mem[4184] = 80'h0010ffabffabffabffab;
mem[4185] = 80'h0010ffabffabffabffab;
mem[4186] = 80'h0010ffabffabffabffab;
mem[4187] = 80'h0010ffabffabffabffab;
mem[4188] = 80'h0010ffabffabffabffab;
mem[4189] = 80'h0010ffabffabffabffab;
mem[4190] = 80'h0010ffabffabffabffab;
mem[4191] = 80'h0010ffabffabffabffab;
mem[4192] = 80'h0010ffabffabffabffab;
mem[4193] = 80'h0010ffabffabffabffab;
mem[4194] = 80'h0010ffabffabffabffab;
mem[4195] = 80'h0010ffabffabffabffab;
mem[4196] = 80'h0010ffabffabffabffab;
mem[4197] = 80'h0010ffabffabffabffab;
mem[4198] = 80'h0010ffabffabffabffab;
mem[4199] = 80'h0010ffabffabffabffab;
mem[4200] = 80'h0010ffabffabffabffab;
mem[4201] = 80'h0010ffabffabffabffab;
mem[4202] = 80'h0010ffabffabffabffab;
mem[4203] = 80'h0010ffabffabffabffab;
mem[4204] = 80'h0010ffabffabffabffab;
mem[4205] = 80'h0010ffabffabffabffab;
mem[4206] = 80'h0010ffabffabffabffab;
mem[4207] = 80'h0010ffabffabffabffab;
mem[4208] = 80'h0010ffabffabffabffab;
mem[4209] = 80'h0010ffabffabffabffab;
mem[4210] = 80'h0010ffabffabffabffab;
mem[4211] = 80'h0010ffabffabffabffab;
mem[4212] = 80'h0010ffabffabffabffab;
mem[4213] = 80'h0010ffabffabffabffab;
mem[4214] = 80'h0010ffabffabffabffab;
mem[4215] = 80'h0010ffabffabffabffab;
mem[4216] = 80'h0010ffabffabffabffab;
mem[4217] = 80'h0010ffabffabffabffab;
mem[4218] = 80'h0010ffabffabffabffab;
mem[4219] = 80'h0010ffabffabffabffab;
mem[4220] = 80'h0010ffabffabffabffab;
mem[4221] = 80'h0010ffabffabffabffab;
mem[4222] = 80'h0010ffabffabffabffab;
mem[4223] = 80'h0010ffabffabffabffab;
mem[4224] = 80'h0010ffabffabffabffab;
mem[4225] = 80'h0010ffabffabffabffab;
mem[4226] = 80'h0010ffabffabffabffab;
mem[4227] = 80'h0010ffabffabffabffab;
mem[4228] = 80'h0010ffabffabffabffab;
mem[4229] = 80'h0010ffabffabffabffab;
mem[4230] = 80'h0010ffabffabffabffab;
mem[4231] = 80'h0010ffabffabffabffab;
mem[4232] = 80'h0010ffabffabffabffab;
mem[4233] = 80'h0010ffabffabffabffab;
mem[4234] = 80'h0010ffabffabffabffab;
mem[4235] = 80'h0010ffabffabffabffab;
mem[4236] = 80'h0010ffabffabffabffab;
mem[4237] = 80'h0010ffabffabffabffab;
mem[4238] = 80'h0010ffabffabffabffab;
mem[4239] = 80'h0010ffabffabffabffab;
mem[4240] = 80'h0010ffabffabffabffab;
mem[4241] = 80'h0010ffabffabffabffab;
mem[4242] = 80'h0010ffabffabffabffab;
mem[4243] = 80'h0010ffabffabffabffab;
mem[4244] = 80'h0010ffabffabffabffab;
mem[4245] = 80'h0010ffabffabffabff3e;
mem[4246] = 80'h001002e2bc59397bf308;
mem[4247] = 80'h00101e64c837a9d0a23c;
mem[4248] = 80'h01176d587489831b1800;
mem[4249] = 80'h10100000010000010010;
mem[4250] = 80'h00109400000208004500;
mem[4251] = 80'h001002bd89c20000fffd;
mem[4252] = 80'h0010ad28c0550102c000;
mem[4253] = 80'h00100001ffabffabffab;
mem[4254] = 80'h0010ffabffabffabffab;
mem[4255] = 80'h0010ffabffabffabffab;
mem[4256] = 80'h0010ffabffabffabffab;
mem[4257] = 80'h0010ffabffabffabffab;
mem[4258] = 80'h0010ffabffabffabffab;
mem[4259] = 80'h0010ffabffabffabffab;
mem[4260] = 80'h0010ffabffabffabffab;
mem[4261] = 80'h0010ffabffabffabffab;
mem[4262] = 80'h0010ffabffabffabffab;
mem[4263] = 80'h0010ffabffabffabffab;
mem[4264] = 80'h0010ffabffabffabffab;
mem[4265] = 80'h0010ffabffabffabffab;
mem[4266] = 80'h0010ffabffabffabffab;
mem[4267] = 80'h0010ffabffabffabffab;
mem[4268] = 80'h0010ffabffabffabffab;
mem[4269] = 80'h0010ffabffabffabffab;
mem[4270] = 80'h0010ffabffabffabffab;
mem[4271] = 80'h0010ffabffabffabffab;
mem[4272] = 80'h0010ffabffabffabffab;
mem[4273] = 80'h0010ffabffabffabffab;
mem[4274] = 80'h0010ffabffabffabffab;
mem[4275] = 80'h0010ffabffabffabffab;
mem[4276] = 80'h0010ffabffabffabffab;
mem[4277] = 80'h0010ffabffabffabffab;
mem[4278] = 80'h0010ffabffabffabffab;
mem[4279] = 80'h0010ffabffabffabffab;
mem[4280] = 80'h0010ffabffabffabffab;
mem[4281] = 80'h0010ffabffabffabffab;
mem[4282] = 80'h0010ffabffabffabffab;
mem[4283] = 80'h0010ffabffabffabffab;
mem[4284] = 80'h0010ffabffabffabffab;
mem[4285] = 80'h0010ffabffabffabffab;
mem[4286] = 80'h0010ffabffabffabffab;
mem[4287] = 80'h0010ffabffabffabffab;
mem[4288] = 80'h0010ffabffabffabffab;
mem[4289] = 80'h0010ffabffabffabffab;
mem[4290] = 80'h0010ffabffabffabffab;
mem[4291] = 80'h0010ffabffabffabffab;
mem[4292] = 80'h0010ffabffabffabffab;
mem[4293] = 80'h0010ffabffabffabffab;
mem[4294] = 80'h0010ffabffabffabffab;
mem[4295] = 80'h0010ffabffabffabffab;
mem[4296] = 80'h0010ffabffabffabffab;
mem[4297] = 80'h0010ffabffabffabffab;
mem[4298] = 80'h0010ffabffabffabffab;
mem[4299] = 80'h0010ffabffabffabffab;
mem[4300] = 80'h0010ffabffabffabffab;
mem[4301] = 80'h0010ffabffabffabffab;
mem[4302] = 80'h0010ffabffabffabffab;
mem[4303] = 80'h0010ffabffabffabffab;
mem[4304] = 80'h0010ffabffabffabffab;
mem[4305] = 80'h0010ffabffabffabffab;
mem[4306] = 80'h0010ffabffabffabffab;
mem[4307] = 80'h0010ffabffabffabffab;
mem[4308] = 80'h0010ffabffabffabffab;
mem[4309] = 80'h0010ffabffabffabffab;
mem[4310] = 80'h0010ffabffabffabffab;
mem[4311] = 80'h0010ffabffabffabffab;
mem[4312] = 80'h0010ffabffabffabffab;
mem[4313] = 80'h0010ffabffabffabffab;
mem[4314] = 80'h0010ffabffabffabffab;
mem[4315] = 80'h0010ffabffabffabffab;
mem[4316] = 80'h0010ffabffabffabffab;
mem[4317] = 80'h0010ffabffabffabffab;
mem[4318] = 80'h0010ffabffabffabffab;
mem[4319] = 80'h0010ffabffabffabffab;
mem[4320] = 80'h0010ffabffabffabffab;
mem[4321] = 80'h0010ffabffabffabffab;
mem[4322] = 80'h0010ffabffabffabffab;
mem[4323] = 80'h0010ffabffabffabffab;
mem[4324] = 80'h0010ffabffabffabffab;
mem[4325] = 80'h0010ffabffabffabffab;
mem[4326] = 80'h0010ffabffabffabffab;
mem[4327] = 80'h0010ffabffabffabffab;
mem[4328] = 80'h0010ffabffabffabffab;
mem[4329] = 80'h0010ffabffabffabffab;
mem[4330] = 80'h0010ffabffabffabffab;
mem[4331] = 80'h0010ffabffabffabffab;
mem[4332] = 80'h0010ffabffabffabffab;
mem[4333] = 80'h0010ffabffabffabffab;
mem[4334] = 80'h0010ffabffabffabffab;
mem[4335] = 80'h0010ffabffabffabff3d;
mem[4336] = 80'h00109080c931b33c3354;
mem[4337] = 80'h001069ecfe29df3f500c;
mem[4338] = 80'h01173e1cea2e26975a00;
mem[4339] = 80'h10100000010000010010;
mem[4340] = 80'h00109400000208004500;
mem[4341] = 80'h0010044d89c30000fffd;
mem[4342] = 80'h0010ab97c0550102c000;
mem[4343] = 80'h00100001ffabffabffab;
mem[4344] = 80'h0010ffabffabffabffab;
mem[4345] = 80'h0010ffabffabffabffab;
mem[4346] = 80'h0010ffabffabffabffab;
mem[4347] = 80'h0010ffabffabffabffab;
mem[4348] = 80'h0010ffabffabffabffab;
mem[4349] = 80'h0010ffabffabffabffab;
mem[4350] = 80'h0010ffabffabffabffab;
mem[4351] = 80'h0010ffabffabffabffab;
mem[4352] = 80'h0010ffabffabffabffab;
mem[4353] = 80'h0010ffabffabffabffab;
mem[4354] = 80'h0010ffabffabffabffab;
mem[4355] = 80'h0010ffabffabffabffab;
mem[4356] = 80'h0010ffabffabffabffab;
mem[4357] = 80'h0010ffabffabffabffab;
mem[4358] = 80'h0010ffabffabffabffab;
mem[4359] = 80'h0010ffabffabffabffab;
mem[4360] = 80'h0010ffabffabffabffab;
mem[4361] = 80'h0010ffabffabffabffab;
mem[4362] = 80'h0010ffabffabffabffab;
mem[4363] = 80'h0010ffabffabffabffab;
mem[4364] = 80'h0010ffabffabffabffab;
mem[4365] = 80'h0010ffabffabffabffab;
mem[4366] = 80'h0010ffabffabffabffab;
mem[4367] = 80'h0010ffabffabffabffab;
mem[4368] = 80'h0010ffabffabffabffab;
mem[4369] = 80'h0010ffabffabffabffab;
mem[4370] = 80'h0010ffabffabffabffab;
mem[4371] = 80'h0010ffabffabffabffab;
mem[4372] = 80'h0010ffabffabffabffab;
mem[4373] = 80'h0010ffabffabffabffab;
mem[4374] = 80'h0010ffabffabffabffab;
mem[4375] = 80'h0010ffabffabffabffab;
mem[4376] = 80'h0010ffabffabffabffab;
mem[4377] = 80'h0010ffabffabffabffab;
mem[4378] = 80'h0010ffabffabffabffab;
mem[4379] = 80'h0010ffabffabffabffab;
mem[4380] = 80'h0010ffabffabffabffab;
mem[4381] = 80'h0010ffabffabffabffab;
mem[4382] = 80'h0010ffabffabffabffab;
mem[4383] = 80'h0010ffabffabffabffab;
mem[4384] = 80'h0010ffabffabffabffab;
mem[4385] = 80'h0010ffabffabffabffab;
mem[4386] = 80'h0010ffabffabffabffab;
mem[4387] = 80'h0010ffabffabffabffab;
mem[4388] = 80'h0010ffabffabffabffab;
mem[4389] = 80'h0010ffabffabffabffab;
mem[4390] = 80'h0010ffabffabffabffab;
mem[4391] = 80'h0010ffabffabffabffab;
mem[4392] = 80'h0010ffabffabffabffab;
mem[4393] = 80'h0010ffabffabffabffab;
mem[4394] = 80'h0010ffabffabffabffab;
mem[4395] = 80'h0010ffabffabffabffab;
mem[4396] = 80'h0010ffabffabffabffab;
mem[4397] = 80'h0010ffabffabffabffab;
mem[4398] = 80'h0010ffabffabffabffab;
mem[4399] = 80'h0010ffabffabffabffab;
mem[4400] = 80'h0010ffabffabffabffab;
mem[4401] = 80'h0010ffabffabffabffab;
mem[4402] = 80'h0010ffabffabffabffab;
mem[4403] = 80'h0010ffabffabffabffab;
mem[4404] = 80'h0010ffabffabffabffab;
mem[4405] = 80'h0010ffabffabffabffab;
mem[4406] = 80'h0010ffabffabffabffab;
mem[4407] = 80'h0010ffabffabffabffab;
mem[4408] = 80'h0010ffabffabffabffab;
mem[4409] = 80'h0010ffabffabffabffab;
mem[4410] = 80'h0010ffabffabffabffab;
mem[4411] = 80'h0010ffabffabffabffab;
mem[4412] = 80'h0010ffabffabffabffab;
mem[4413] = 80'h0010ffabffabffabffab;
mem[4414] = 80'h0010ffabffabffabffab;
mem[4415] = 80'h0010ffabffabffabffab;
mem[4416] = 80'h0010ffabffabffabffab;
mem[4417] = 80'h0010ffabffabffabffab;
mem[4418] = 80'h0010ffabffabffabffab;
mem[4419] = 80'h0010ffabffabffabffab;
mem[4420] = 80'h0010ffabffabffabffab;
mem[4421] = 80'h0010ffabffabffabffab;
mem[4422] = 80'h0010ffabffabffabffab;
mem[4423] = 80'h0010ffabffabffabffab;
mem[4424] = 80'h0010ffabffabffabffab;
mem[4425] = 80'h0010ffabffabffabffab;
mem[4426] = 80'h0010ffabffabffabffab;
mem[4427] = 80'h0010ffabffabffabffab;
mem[4428] = 80'h0010ffabffabffabffab;
mem[4429] = 80'h0010ffabffabffabffab;
mem[4430] = 80'h0010ffabffabffabffab;
mem[4431] = 80'h0010ffabffabffabffab;
mem[4432] = 80'h0010ffabffabffabffab;
mem[4433] = 80'h0010ffabffabffabffab;
mem[4434] = 80'h0010ffabffabffabffab;
mem[4435] = 80'h0010ffabffabffabffab;
mem[4436] = 80'h0010ffabffabffabffab;
mem[4437] = 80'h0010ffabffabffabffab;
mem[4438] = 80'h0010ffabffabffabffab;
mem[4439] = 80'h0010ffabffabffabffab;
mem[4440] = 80'h0010ffabffabffabffab;
mem[4441] = 80'h0010ffabffabffabffab;
mem[4442] = 80'h0010ffabffabffabffab;
mem[4443] = 80'h0010ffabffabffabffab;
mem[4444] = 80'h0010ffabffabffabffab;
mem[4445] = 80'h0010ffabffabffabffab;
mem[4446] = 80'h0010ffabffabffabffab;
mem[4447] = 80'h0010ffabffabffabffab;
mem[4448] = 80'h0010ffabffabffabffab;
mem[4449] = 80'h0010ffabffabffabffab;
mem[4450] = 80'h0010ffabffabffabffab;
mem[4451] = 80'h0010ffabffabffabffab;
mem[4452] = 80'h0010ffabffabffabffab;
mem[4453] = 80'h0010ffabffabffabffab;
mem[4454] = 80'h0010ffabffabffabffab;
mem[4455] = 80'h0010ffabffabffabffab;
mem[4456] = 80'h0010ffabffabffabffab;
mem[4457] = 80'h0010ffabffabffabffab;
mem[4458] = 80'h0010ffabffabffabffab;
mem[4459] = 80'h0010ffabffabffabffab;
mem[4460] = 80'h0010ffabffabffabffab;
mem[4461] = 80'h0010ffabffabffabffab;
mem[4462] = 80'h0010ffabffabffabffab;
mem[4463] = 80'h0010ffabffabffabffab;
mem[4464] = 80'h0010ffabffabffabffab;
mem[4465] = 80'h0010ffabffabffabffab;
mem[4466] = 80'h0010ffabffabffabffab;
mem[4467] = 80'h0010ffabffabffabffab;
mem[4468] = 80'h0010ffabffabffabffab;
mem[4469] = 80'h0010ffabffabffabffab;
mem[4470] = 80'h0010ffabffabffabffab;
mem[4471] = 80'h0010ffabffabffabffab;
mem[4472] = 80'h0010ffabffabffabffab;
mem[4473] = 80'h0010ffabffabffabffab;
mem[4474] = 80'h0010ffabffabffabffab;
mem[4475] = 80'h0010ffabffabffabff3c;
mem[4476] = 80'h0010e15ee5e9cafe8c9f;
mem[4477] = 80'h0010bb6b13dc0e7601fd;
mem[4478] = 80'h011790217151192e5500;
mem[4479] = 80'h10100000010000010010;
mem[4480] = 80'h00109400000208004500;
mem[4481] = 80'h0010023d89c40000fffd;
mem[4482] = 80'h0010ada6c0550102c000;
mem[4483] = 80'h00100001ffabffabffab;
mem[4484] = 80'h0010ffabffabffabffab;
mem[4485] = 80'h0010ffabffabffabffab;
mem[4486] = 80'h0010ffabffabffabffab;
mem[4487] = 80'h0010ffabffabffabffab;
mem[4488] = 80'h0010ffabffabffabffab;
mem[4489] = 80'h0010ffabffabffabffab;
mem[4490] = 80'h0010ffabffabffabffab;
mem[4491] = 80'h0010ffabffabffabffab;
mem[4492] = 80'h0010ffabffabffabffab;
mem[4493] = 80'h0010ffabffabffabffab;
mem[4494] = 80'h0010ffabffabffabffab;
mem[4495] = 80'h0010ffabffabffabffab;
mem[4496] = 80'h0010ffabffabffabffab;
mem[4497] = 80'h0010ffabffabffabffab;
mem[4498] = 80'h0010ffabffabffabffab;
mem[4499] = 80'h0010ffabffabffabffab;
mem[4500] = 80'h0010ffabffabffabffab;
mem[4501] = 80'h0010ffabffabffabffab;
mem[4502] = 80'h0010ffabffabffabffab;
mem[4503] = 80'h0010ffabffabffabffab;
mem[4504] = 80'h0010ffabffabffabffab;
mem[4505] = 80'h0010ffabffabffabffab;
mem[4506] = 80'h0010ffabffabffabffab;
mem[4507] = 80'h0010ffabffabffabffab;
mem[4508] = 80'h0010ffabffabffabffab;
mem[4509] = 80'h0010ffabffabffabffab;
mem[4510] = 80'h0010ffabffabffabffab;
mem[4511] = 80'h0010ffabffabffabffab;
mem[4512] = 80'h0010ffabffabffabffab;
mem[4513] = 80'h0010ffabffabffabffab;
mem[4514] = 80'h0010ffabffabffabffab;
mem[4515] = 80'h0010ffabffabffabffab;
mem[4516] = 80'h0010ffabffabffabffab;
mem[4517] = 80'h0010ffabffabffabffab;
mem[4518] = 80'h0010ffabffabffabffab;
mem[4519] = 80'h0010ffabffabffabffab;
mem[4520] = 80'h0010ffabffabffabffab;
mem[4521] = 80'h0010ffabffabffabffab;
mem[4522] = 80'h0010ffabffabffabffab;
mem[4523] = 80'h0010ffabffabffabffab;
mem[4524] = 80'h0010ffabffabffabffab;
mem[4525] = 80'h0010ffabffabffabffab;
mem[4526] = 80'h0010ffabffabffabffab;
mem[4527] = 80'h0010ffabffabffabffab;
mem[4528] = 80'h0010ffabffabffabffab;
mem[4529] = 80'h0010ffabffabffabffab;
mem[4530] = 80'h0010ffabffabffabffab;
mem[4531] = 80'h0010ffabffabffabffab;
mem[4532] = 80'h0010ffabffabffabffab;
mem[4533] = 80'h0010ffabffabffabffab;
mem[4534] = 80'h0010ffabffabffabffab;
mem[4535] = 80'h0010ffabffabffabffab;
mem[4536] = 80'h0010ffabffabffabffab;
mem[4537] = 80'h0010ffabffabffabffab;
mem[4538] = 80'h0010ffabffabffabffab;
mem[4539] = 80'h0010ffabffabffabffab;
mem[4540] = 80'h0010ffabffabffabffab;
mem[4541] = 80'h0010ffabffabffabffab;
mem[4542] = 80'h0010ffabffabffabffab;
mem[4543] = 80'h0010ffabffabffabffab;
mem[4544] = 80'h0010ffabffabffabffab;
mem[4545] = 80'h0010ffabffabffabffab;
mem[4546] = 80'h0010ffabffabffabffab;
mem[4547] = 80'h0010ffabffabffabffab;
mem[4548] = 80'h0010ffabffabffabffab;
mem[4549] = 80'h0010ffabffabffabff3b;
mem[4550] = 80'h0010c59a0f38de710c27;
mem[4551] = 80'h0010547a7fe0ecbce418;
mem[4552] = 80'h011700289ba2b4957900;
mem[4553] = 80'h10100000010000010010;
mem[4554] = 80'h00109400000208004500;
mem[4555] = 80'h0010040d89c50000fffd;
mem[4556] = 80'h0010abd5c0550102c000;
mem[4557] = 80'h00100001ffabffabffab;
mem[4558] = 80'h0010ffabffabffabffab;
mem[4559] = 80'h0010ffabffabffabffab;
mem[4560] = 80'h0010ffabffabffabffab;
mem[4561] = 80'h0010ffabffabffabffab;
mem[4562] = 80'h0010ffabffabffabffab;
mem[4563] = 80'h0010ffabffabffabffab;
mem[4564] = 80'h0010ffabffabffabffab;
mem[4565] = 80'h0010ffabffabffabffab;
mem[4566] = 80'h0010ffabffabffabffab;
mem[4567] = 80'h0010ffabffabffabffab;
mem[4568] = 80'h0010ffabffabffabffab;
mem[4569] = 80'h0010ffabffabffabffab;
mem[4570] = 80'h0010ffabffabffabffab;
mem[4571] = 80'h0010ffabffabffabffab;
mem[4572] = 80'h0010ffabffabffabffab;
mem[4573] = 80'h0010ffabffabffabffab;
mem[4574] = 80'h0010ffabffabffabffab;
mem[4575] = 80'h0010ffabffabffabffab;
mem[4576] = 80'h0010ffabffabffabffab;
mem[4577] = 80'h0010ffabffabffabffab;
mem[4578] = 80'h0010ffabffabffabffab;
mem[4579] = 80'h0010ffabffabffabffab;
mem[4580] = 80'h0010ffabffabffabffab;
mem[4581] = 80'h0010ffabffabffabffab;
mem[4582] = 80'h0010ffabffabffabffab;
mem[4583] = 80'h0010ffabffabffabffab;
mem[4584] = 80'h0010ffabffabffabffab;
mem[4585] = 80'h0010ffabffabffabffab;
mem[4586] = 80'h0010ffabffabffabffab;
mem[4587] = 80'h0010ffabffabffabffab;
mem[4588] = 80'h0010ffabffabffabffab;
mem[4589] = 80'h0010ffabffabffabffab;
mem[4590] = 80'h0010ffabffabffabffab;
mem[4591] = 80'h0010ffabffabffabffab;
mem[4592] = 80'h0010ffabffabffabffab;
mem[4593] = 80'h0010ffabffabffabffab;
mem[4594] = 80'h0010ffabffabffabffab;
mem[4595] = 80'h0010ffabffabffabffab;
mem[4596] = 80'h0010ffabffabffabffab;
mem[4597] = 80'h0010ffabffabffabffab;
mem[4598] = 80'h0010ffabffabffabffab;
mem[4599] = 80'h0010ffabffabffabffab;
mem[4600] = 80'h0010ffabffabffabffab;
mem[4601] = 80'h0010ffabffabffabffab;
mem[4602] = 80'h0010ffabffabffabffab;
mem[4603] = 80'h0010ffabffabffabffab;
mem[4604] = 80'h0010ffabffabffabffab;
mem[4605] = 80'h0010ffabffabffabffab;
mem[4606] = 80'h0010ffabffabffabffab;
mem[4607] = 80'h0010ffabffabffabffab;
mem[4608] = 80'h0010ffabffabffabffab;
mem[4609] = 80'h0010ffabffabffabffab;
mem[4610] = 80'h0010ffabffabffabffab;
mem[4611] = 80'h0010ffabffabffabffab;
mem[4612] = 80'h0010ffabffabffabffab;
mem[4613] = 80'h0010ffabffabffabffab;
mem[4614] = 80'h0010ffabffabffabffab;
mem[4615] = 80'h0010ffabffabffabffab;
mem[4616] = 80'h0010ffabffabffabffab;
mem[4617] = 80'h0010ffabffabffabffab;
mem[4618] = 80'h0010ffabffabffabffab;
mem[4619] = 80'h0010ffabffabffabffab;
mem[4620] = 80'h0010ffabffabffabffab;
mem[4621] = 80'h0010ffabffabffabffab;
mem[4622] = 80'h0010ffabffabffabffab;
mem[4623] = 80'h0010ffabffabffabffab;
mem[4624] = 80'h0010ffabffabffabffab;
mem[4625] = 80'h0010ffabffabffabffab;
mem[4626] = 80'h0010ffabffabffabffab;
mem[4627] = 80'h0010ffabffabffabffab;
mem[4628] = 80'h0010ffabffabffabffab;
mem[4629] = 80'h0010ffabffabffabffab;
mem[4630] = 80'h0010ffabffabffabffab;
mem[4631] = 80'h0010ffabffabffabffab;
mem[4632] = 80'h0010ffabffabffabffab;
mem[4633] = 80'h0010ffabffabffabffab;
mem[4634] = 80'h0010ffabffabffabffab;
mem[4635] = 80'h0010ffabffabffabffab;
mem[4636] = 80'h0010ffabffabffabffab;
mem[4637] = 80'h0010ffabffabffabffab;
mem[4638] = 80'h0010ffabffabffabffab;
mem[4639] = 80'h0010ffabffabffabffab;
mem[4640] = 80'h0010ffabffabffabffab;
mem[4641] = 80'h0010ffabffabffabffab;
mem[4642] = 80'h0010ffabffabffabffab;
mem[4643] = 80'h0010ffabffabffabffab;
mem[4644] = 80'h0010ffabffabffabffab;
mem[4645] = 80'h0010ffabffabffabffab;
mem[4646] = 80'h0010ffabffabffabffab;
mem[4647] = 80'h0010ffabffabffabffab;
mem[4648] = 80'h0010ffabffabffabffab;
mem[4649] = 80'h0010ffabffabffabffab;
mem[4650] = 80'h0010ffabffabffabffab;
mem[4651] = 80'h0010ffabffabffabffab;
mem[4652] = 80'h0010ffabffabffabffab;
mem[4653] = 80'h0010ffabffabffabffab;
mem[4654] = 80'h0010ffabffabffabffab;
mem[4655] = 80'h0010ffabffabffabffab;
mem[4656] = 80'h0010ffabffabffabffab;
mem[4657] = 80'h0010ffabffabffabffab;
mem[4658] = 80'h0010ffabffabffabffab;
mem[4659] = 80'h0010ffabffabffabffab;
mem[4660] = 80'h0010ffabffabffabffab;
mem[4661] = 80'h0010ffabffabffabffab;
mem[4662] = 80'h0010ffabffabffabffab;
mem[4663] = 80'h0010ffabffabffabffab;
mem[4664] = 80'h0010ffabffabffabffab;
mem[4665] = 80'h0010ffabffabffabffab;
mem[4666] = 80'h0010ffabffabffabffab;
mem[4667] = 80'h0010ffabffabffabffab;
mem[4668] = 80'h0010ffabffabffabffab;
mem[4669] = 80'h0010ffabffabffabffab;
mem[4670] = 80'h0010ffabffabffabffab;
mem[4671] = 80'h0010ffabffabffabffab;
mem[4672] = 80'h0010ffabffabffabffab;
mem[4673] = 80'h0010ffabffabffabffab;
mem[4674] = 80'h0010ffabffabffabffab;
mem[4675] = 80'h0010ffabffabffabffab;
mem[4676] = 80'h0010ffabffabffabffab;
mem[4677] = 80'h0010ffabffabffabffab;
mem[4678] = 80'h0010ffabffabffabffab;
mem[4679] = 80'h0010ffabffabffabffab;
mem[4680] = 80'h0010ffabffabffabffab;
mem[4681] = 80'h0010ffabffabffabff3a;
mem[4682] = 80'h0010b44423e0a7b3b3ec;
mem[4683] = 80'h001086fd92153d1cb543;
mem[4684] = 80'h0117848d3c37b4e3b500;
mem[4685] = 80'h10100000010000010010;
mem[4686] = 80'h00109400000208004500;
mem[4687] = 80'h0010021f89c60000fffd;
mem[4688] = 80'h0010adc2c0550102c000;
mem[4689] = 80'h00100001ffabffabffab;
mem[4690] = 80'h0010ffabffabffabffab;
mem[4691] = 80'h0010ffabffabffabffab;
mem[4692] = 80'h0010ffabffabffabffab;
mem[4693] = 80'h0010ffabffabffabffab;
mem[4694] = 80'h0010ffabffabffabffab;
mem[4695] = 80'h0010ffabffabffabffab;
mem[4696] = 80'h0010ffabffabffabffab;
mem[4697] = 80'h0010ffabffabffabffab;
mem[4698] = 80'h0010ffabffabffabffab;
mem[4699] = 80'h0010ffabffabffabffab;
mem[4700] = 80'h0010ffabffabffabffab;
mem[4701] = 80'h0010ffabffabffabffab;
mem[4702] = 80'h0010ffabffabffabffab;
mem[4703] = 80'h0010ffabffabffabffab;
mem[4704] = 80'h0010ffabffabffabffab;
mem[4705] = 80'h0010ffabffabffabffab;
mem[4706] = 80'h0010ffabffabffabffab;
mem[4707] = 80'h0010ffabffabffabffab;
mem[4708] = 80'h0010ffabffabffabffab;
mem[4709] = 80'h0010ffabffabffabffab;
mem[4710] = 80'h0010ffabffabffabffab;
mem[4711] = 80'h0010ffabffabffabffab;
mem[4712] = 80'h0010ffabffabffabffab;
mem[4713] = 80'h0010ffabffabffabffab;
mem[4714] = 80'h0010ffabffabffabffab;
mem[4715] = 80'h0010ffabffabffabffab;
mem[4716] = 80'h0010ffabffabffabffab;
mem[4717] = 80'h0010ffabffabffabffab;
mem[4718] = 80'h0010ffabffabffabffab;
mem[4719] = 80'h0010ffabffabffabffab;
mem[4720] = 80'h0010ffabffabffabffab;
mem[4721] = 80'h0010ffabffabffabffab;
mem[4722] = 80'h0010ffabffabffabffab;
mem[4723] = 80'h0010ffabffabffabffab;
mem[4724] = 80'h0010ffabffabffabffab;
mem[4725] = 80'h0010ffabffabffabffab;
mem[4726] = 80'h0010ffabffabffabffab;
mem[4727] = 80'h0010ffabffabffabffab;
mem[4728] = 80'h0010ffabffabffabffab;
mem[4729] = 80'h0010ffabffabffabffab;
mem[4730] = 80'h0010ffabffabffabffab;
mem[4731] = 80'h0010ffabffabffabffab;
mem[4732] = 80'h0010ffabffabffabffab;
mem[4733] = 80'h0010ffabffabffabffab;
mem[4734] = 80'h0010ffabffabffabffab;
mem[4735] = 80'h0010ffabffabffabffab;
mem[4736] = 80'h0010ffabffabffabffab;
mem[4737] = 80'h0010ffabffabffabffab;
mem[4738] = 80'h0010ffabffabffabffab;
mem[4739] = 80'h0010ffabffabffabffab;
mem[4740] = 80'h0010ffabffabffabffab;
mem[4741] = 80'h0010ffabffabffabffab;
mem[4742] = 80'h0010ffabffabffabffab;
mem[4743] = 80'h0010ffabffabffabffab;
mem[4744] = 80'h0010ffabffabffabffab;
mem[4745] = 80'h0010ffabffabffabffab;
mem[4746] = 80'h0010ffabffabffabffab;
mem[4747] = 80'h0010ffabffabffabffab;
mem[4748] = 80'h0010ffabffabffabffab;
mem[4749] = 80'h0010ffabffabffabffab;
mem[4750] = 80'h0010ffabffabffabffab;
mem[4751] = 80'h0010ffabffabffabffab;
mem[4752] = 80'h0010ff39262656882df4;
mem[4753] = 80'h001073b0f175a40b425a;
mem[4754] = 80'h0010474aa04d2288b12a;
mem[4755] = 80'h0111a400000000000000;
mem[4756] = 80'h10100000010000010010;
mem[4757] = 80'h00109400000208004500;
mem[4758] = 80'h001003ff89c70000fffd;
mem[4759] = 80'h0010abe1c0550102c000;
mem[4760] = 80'h00100001ffabffabffab;
mem[4761] = 80'h0010ffabffabffabffab;
mem[4762] = 80'h0010ffabffabffabffab;
mem[4763] = 80'h0010ffabffabffabffab;
mem[4764] = 80'h0010ffabffabffabffab;
mem[4765] = 80'h0010ffabffabffabffab;
mem[4766] = 80'h0010ffabffabffabffab;
mem[4767] = 80'h0010ffabffabffabffab;
mem[4768] = 80'h0010ffabffabffabffab;
mem[4769] = 80'h0010ffabffabffabffab;
mem[4770] = 80'h0010ffabffabffabffab;
mem[4771] = 80'h0010ffabffabffabffab;
mem[4772] = 80'h0010ffabffabffabffab;
mem[4773] = 80'h0010ffabffabffabffab;
mem[4774] = 80'h0010ffabffabffabffab;
mem[4775] = 80'h0010ffabffabffabffab;
mem[4776] = 80'h0010ffabffabffabffab;
mem[4777] = 80'h0010ffabffabffabffab;
mem[4778] = 80'h0010ffabffabffabffab;
mem[4779] = 80'h0010ffabffabffabffab;
mem[4780] = 80'h0010ffabffabffabffab;
mem[4781] = 80'h0010ffabffabffabffab;
mem[4782] = 80'h0010ffabffabffabffab;
mem[4783] = 80'h0010ffabffabffabffab;
mem[4784] = 80'h0010ffabffabffabffab;
mem[4785] = 80'h0010ffabffabffabffab;
mem[4786] = 80'h0010ffabffabffabffab;
mem[4787] = 80'h0010ffabffabffabffab;
mem[4788] = 80'h0010ffabffabffabffab;
mem[4789] = 80'h0010ffabffabffabffab;
mem[4790] = 80'h0010ffabffabffabffab;
mem[4791] = 80'h0010ffabffabffabffab;
mem[4792] = 80'h0010ffabffabffabffab;
mem[4793] = 80'h0010ffabffabffabffab;
mem[4794] = 80'h0010ffabffabffabffab;
mem[4795] = 80'h0010ffabffabffabffab;
mem[4796] = 80'h0010ffabffabffabffab;
mem[4797] = 80'h0010ffabffabffabffab;
mem[4798] = 80'h0010ffabffabffabffab;
mem[4799] = 80'h0010ffabffabffabffab;
mem[4800] = 80'h0010ffabffabffabffab;
mem[4801] = 80'h0010ffabffabffabffab;
mem[4802] = 80'h0010ffabffabffabffab;
mem[4803] = 80'h0010ffabffabffabffab;
mem[4804] = 80'h0010ffabffabffabffab;
mem[4805] = 80'h0010ffabffabffabffab;
mem[4806] = 80'h0010ffabffabffabffab;
mem[4807] = 80'h0010ffabffabffabffab;
mem[4808] = 80'h0010ffabffabffabffab;
mem[4809] = 80'h0010ffabffabffabffab;
mem[4810] = 80'h0010ffabffabffabffab;
mem[4811] = 80'h0010ffabffabffabffab;
mem[4812] = 80'h0010ffabffabffabffab;
mem[4813] = 80'h0010ffabffabffabffab;
mem[4814] = 80'h0010ffabffabffabffab;
mem[4815] = 80'h0010ffabffabffabffab;
mem[4816] = 80'h0010ffabffabffabffab;
mem[4817] = 80'h0010ffabffabffabffab;
mem[4818] = 80'h0010ffabffabffabffab;
mem[4819] = 80'h0010ffabffabffabffab;
mem[4820] = 80'h0010ffabffabffabffab;
mem[4821] = 80'h0010ffabffabffabffab;
mem[4822] = 80'h0010ffabffabffabffab;
mem[4823] = 80'h0010ffabffabffabffab;
mem[4824] = 80'h0010ffabffabffabffab;
mem[4825] = 80'h0010ffabffabffabffab;
mem[4826] = 80'h0010ffabffabffabffab;
mem[4827] = 80'h0010ffabffabffabffab;
mem[4828] = 80'h0010ffabffabffabffab;
mem[4829] = 80'h0010ffabffabffabffab;
mem[4830] = 80'h0010ffabffabffabffab;
mem[4831] = 80'h0010ffabffabffabffab;
mem[4832] = 80'h0010ffabffabffabffab;
mem[4833] = 80'h0010ffabffabffabffab;
mem[4834] = 80'h0010ffabffabffabffab;
mem[4835] = 80'h0010ffabffabffabffab;
mem[4836] = 80'h0010ffabffabffabffab;
mem[4837] = 80'h0010ffabffabffabffab;
mem[4838] = 80'h0010ffabffabffabffab;
mem[4839] = 80'h0010ffabffabffabffab;
mem[4840] = 80'h0010ffabffabffabffab;
mem[4841] = 80'h0010ffabffabffabffab;
mem[4842] = 80'h0010ffabffabffabffab;
mem[4843] = 80'h0010ffabffabffabffab;
mem[4844] = 80'h0010ffabffabffabffab;
mem[4845] = 80'h0010ffabffabffabffab;
mem[4846] = 80'h0010ffabffabffabffab;
mem[4847] = 80'h0010ffabffabffabffab;
mem[4848] = 80'h0010ffabffabffabffab;
mem[4849] = 80'h0010ffabffabffabffab;
mem[4850] = 80'h0010ffabffabffabffab;
mem[4851] = 80'h0010ffabffabffabffab;
mem[4852] = 80'h0010ffabffabffabffab;
mem[4853] = 80'h0010ffabffabffabffab;
mem[4854] = 80'h0010ffabffabffabffab;
mem[4855] = 80'h0010ffabffabffabffab;
mem[4856] = 80'h0010ffabffabffabffab;
mem[4857] = 80'h0010ffabffabffabffab;
mem[4858] = 80'h0010ffabffabffabffab;
mem[4859] = 80'h0010ffabffabffabffab;
mem[4860] = 80'h0010ffabffabffabffab;
mem[4861] = 80'h0010ffabffabffabffab;
mem[4862] = 80'h0010ffabffabffabffab;
mem[4863] = 80'h0010ffabffabffabffab;
mem[4864] = 80'h0010ffabffabffabffab;
mem[4865] = 80'h0010ffabffabffabffab;
mem[4866] = 80'h0010ffabffabffabffab;
mem[4867] = 80'h0010ffabffabffabffab;
mem[4868] = 80'h0010ffabffabffabffab;
mem[4869] = 80'h0010ffabffabffabffab;
mem[4870] = 80'h0010ffabffabffabffab;
mem[4871] = 80'h0010ffabffabffabffab;
mem[4872] = 80'h0010ffabffabffabffab;
mem[4873] = 80'h0010ffabffabffabffab;
mem[4874] = 80'h0010ffabffabffabffab;
mem[4875] = 80'h0010ffabffabffabffab;
mem[4876] = 80'h0010ffabffabffabffab;
mem[4877] = 80'h0010ffabffabffabffab;
mem[4878] = 80'h0010ffabffabffabffab;
mem[4879] = 80'h0010ffabffabffabffab;
mem[4880] = 80'h0010ffabffabffabffab;
mem[4881] = 80'h0010ffabffabffabffab;
mem[4882] = 80'h0010ffabffabffabffab;
mem[4883] = 80'h0010ff3857f87a505436;
mem[4884] = 80'h0010cc7b23f249fe93fa;
mem[4885] = 80'h0010161124d0d000946b;
mem[4886] = 80'h0111b500000000000000;
mem[4887] = 80'h00000000000000000000;
mem[4888] = 80'h00000000000000000000;
mem[4889] = 80'h00000000000000000000;
mem[4890] = 80'h00000000000000000000;
mem[4891] = 80'h00000000000000000000;
mem[4892] = 80'h10100000010000010010;
mem[4893] = 80'h00109400000208004500;
mem[4894] = 80'h001004ec89c80000fffd;
mem[4895] = 80'h0010aaf3c0550102c000;
mem[4896] = 80'h00100001ffabffabffab;
mem[4897] = 80'h0010ffabffabffabffab;
mem[4898] = 80'h0010ffabffabffabffab;
mem[4899] = 80'h0010ffabffabffabffab;
mem[4900] = 80'h0010ffabffabffabffab;
mem[4901] = 80'h0010ffabffabffabffab;
mem[4902] = 80'h0010ffabffabffabffab;
mem[4903] = 80'h0010ffabffabffabffab;
mem[4904] = 80'h0010ffabffabffabffab;
mem[4905] = 80'h0010ffabffabffabffab;
mem[4906] = 80'h0010ffabffabffabffab;
mem[4907] = 80'h0010ffabffabffabffab;
mem[4908] = 80'h0010ffabffabffabffab;
mem[4909] = 80'h0010ffabffabffabffab;
mem[4910] = 80'h0010ffabffabffabffab;
mem[4911] = 80'h0010ffabffabffabffab;
mem[4912] = 80'h0010ffabffabffabffab;
mem[4913] = 80'h0010ffabffabffabffab;
mem[4914] = 80'h0010ffabffabffabffab;
mem[4915] = 80'h0010ffabffabffabffab;
mem[4916] = 80'h0010ffabffabffabffab;
mem[4917] = 80'h0010ffabffabffabffab;
mem[4918] = 80'h0010ffabffabffabffab;
mem[4919] = 80'h0010ffabffabffabffab;
mem[4920] = 80'h0010ffabffabffabffab;
mem[4921] = 80'h0010ffabffabffabffab;
mem[4922] = 80'h0010ffabffabffabffab;
mem[4923] = 80'h0010ffabffabffabffab;
mem[4924] = 80'h0010ffabffabffabffab;
mem[4925] = 80'h0010ffabffabffabffab;
mem[4926] = 80'h0010ffabffabffabffab;
mem[4927] = 80'h0010ffabffabffabffab;
mem[4928] = 80'h0010ffabffabffabffab;
mem[4929] = 80'h0010ffabffabffabffab;
mem[4930] = 80'h0010ffabffabffabffab;
mem[4931] = 80'h0010ffabffabffabffab;
mem[4932] = 80'h0010ffabffabffabffab;
mem[4933] = 80'h0010ffabffabffabffab;
mem[4934] = 80'h0010ffabffabffabffab;
mem[4935] = 80'h0010ffabffabffabffab;
mem[4936] = 80'h0010ffabffabffabffab;
mem[4937] = 80'h0010ffabffabffabffab;
mem[4938] = 80'h0010ffabffabffabffab;
mem[4939] = 80'h0010ffabffabffabffab;
mem[4940] = 80'h0010ffabffabffabffab;
mem[4941] = 80'h0010ffabffabffabffab;
mem[4942] = 80'h0010ffabffabffabffab;
mem[4943] = 80'h0010ffabffabffabffab;
mem[4944] = 80'h0010ffabffabffabffab;
mem[4945] = 80'h0010ffabffabffabffab;
mem[4946] = 80'h0010ffabffabffabffab;
mem[4947] = 80'h0010ffabffabffabffab;
mem[4948] = 80'h0010ffabffabffabffab;
mem[4949] = 80'h0010ffabffabffabffab;
mem[4950] = 80'h0010ffabffabffabffab;
mem[4951] = 80'h0010ffabffabffabffab;
mem[4952] = 80'h0010ffabffabffabffab;
mem[4953] = 80'h0010ffabffabffabffab;
mem[4954] = 80'h0010ffabffabffabffab;
mem[4955] = 80'h0010ffabffabffabffab;
mem[4956] = 80'h0010ffabffabffabffab;
mem[4957] = 80'h0010ffabffabffabffab;
mem[4958] = 80'h0010ffabffabffabffab;
mem[4959] = 80'h0010ffabffabffabffab;
mem[4960] = 80'h0010ffabffabffabffab;
mem[4961] = 80'h0010ffabffabffabffab;
mem[4962] = 80'h0010ffabffabffabffab;
mem[4963] = 80'h0010ffabffabffabffab;
mem[4964] = 80'h0010ffabffabffabffab;
mem[4965] = 80'h0010ffabffabffabffab;
mem[4966] = 80'h0010ffabffabffabffab;
mem[4967] = 80'h0010ffabffabffabffab;
mem[4968] = 80'h0010ffabffabffabffab;
mem[4969] = 80'h0010ffabffabffabffab;
mem[4970] = 80'h0010ffabffabffabffab;
mem[4971] = 80'h0010ffabffabffabffab;
mem[4972] = 80'h0010ffabffabffabffab;
mem[4973] = 80'h0010ffabffabffabffab;
mem[4974] = 80'h0010ffabffabffabffab;
mem[4975] = 80'h0010ffabffabffabffab;
mem[4976] = 80'h0010ffabffabffabffab;
mem[4977] = 80'h0010ffabffabffabffab;
mem[4978] = 80'h0010ffabffabffabffab;
mem[4979] = 80'h0010ffabffabffabffab;
mem[4980] = 80'h0010ffabffabffabffab;
mem[4981] = 80'h0010ffabffabffabffab;
mem[4982] = 80'h0010ffabffabffabffab;
mem[4983] = 80'h0010ffabffabffabffab;
mem[4984] = 80'h0010ffabffabffabffab;
mem[4985] = 80'h0010ffabffabffabffab;
mem[4986] = 80'h0010ffabffabffabffab;
mem[4987] = 80'h0010ffabffabffabffab;
mem[4988] = 80'h0010ffabffabffabffab;
mem[4989] = 80'h0010ffabffabffabffab;
mem[4990] = 80'h0010ffabffabffabffab;
mem[4991] = 80'h0010ffabffabffabffab;
mem[4992] = 80'h0010ffabffabffabffab;
mem[4993] = 80'h0010ffabffabffabffab;
mem[4994] = 80'h0010ffabffabffabffab;
mem[4995] = 80'h0010ffabffabffabffab;
mem[4996] = 80'h0010ffabffabffabffab;
mem[4997] = 80'h0010ffabffabffabffab;
mem[4998] = 80'h0010ffabffabffabffab;
mem[4999] = 80'h0010ffabffabffabffab;
mem[5000] = 80'h0010ffabffabffabffab;
mem[5001] = 80'h0010ffabffabffabffab;
mem[5002] = 80'h0010ffabffabffabffab;
mem[5003] = 80'h0010ffabffabffabffab;
mem[5004] = 80'h0010ffabffabffabffab;
mem[5005] = 80'h0010ffabffabffabffab;
mem[5006] = 80'h0010ffabffabffabffab;
mem[5007] = 80'h0010ffabffabffabffab;
mem[5008] = 80'h0010ffabffabffabffab;
mem[5009] = 80'h0010ffabffabffabffab;
mem[5010] = 80'h0010ffabffabffabffab;
mem[5011] = 80'h0010ffabffabffabffab;
mem[5012] = 80'h0010ffabffabffabffab;
mem[5013] = 80'h0010ffabffabffabffab;
mem[5014] = 80'h0010ffabffabffabffab;
mem[5015] = 80'h0010ffabffabffabffab;
mem[5016] = 80'h0010ffabffabffabffab;
mem[5017] = 80'h0010ffabffabffabffab;
mem[5018] = 80'h0010ffabffabffabffab;
mem[5019] = 80'h0010ffabffabffabffab;
mem[5020] = 80'h0010ffabffabffabffab;
mem[5021] = 80'h0010ffabffabffabffab;
mem[5022] = 80'h0010ffabffabffabffab;
mem[5023] = 80'h0010ffabffabffabffab;
mem[5024] = 80'h0010ffabffabffabffab;
mem[5025] = 80'h0010ffabffabffabffab;
mem[5026] = 80'h0010ffabffabffabffab;
mem[5027] = 80'h0010ffabffabffabffab;
mem[5028] = 80'h0010ffabffabffabffab;
mem[5029] = 80'h0010ffabffabffabffab;
mem[5030] = 80'h0010ffabffabffabffab;
mem[5031] = 80'h0010ffabffabffabffab;
mem[5032] = 80'h0010ffabffabffabffab;
mem[5033] = 80'h0010ffabffabffabffab;
mem[5034] = 80'h0010ffabffabffabffab;
mem[5035] = 80'h0010ffabffabffabffab;
mem[5036] = 80'h0010ffabffabffabffab;
mem[5037] = 80'h0010ffabffabffabffab;
mem[5038] = 80'h0010ffabffabffabffab;
mem[5039] = 80'h0010ffabffabffabffab;
mem[5040] = 80'h0010ffabffabffabffab;
mem[5041] = 80'h0010ffabffabffabffab;
mem[5042] = 80'h0010ffabffabffabffab;
mem[5043] = 80'h0010ffabffabffabffab;
mem[5044] = 80'h0010ffabffabffabffab;
mem[5045] = 80'h0010ffabffabffabffab;
mem[5046] = 80'h0010ffabffabffabffab;
mem[5047] = 80'h0010ffabffabffabffab;
mem[5048] = 80'h0010ffabffabffab376f;
mem[5049] = 80'h0010af832a04eb72c12f;
mem[5050] = 80'h0010577c7282f58c802e;
mem[5051] = 80'h011602ac525fb9d50000;
mem[5052] = 80'h10100000010000010010;
mem[5053] = 80'h00109400000208004500;
mem[5054] = 80'h0010028b89c90000fffd;
mem[5055] = 80'h0010ad53c0550102c000;
mem[5056] = 80'h00100001ffabffabffab;
mem[5057] = 80'h0010ffabffabffabffab;
mem[5058] = 80'h0010ffabffabffabffab;
mem[5059] = 80'h0010ffabffabffabffab;
mem[5060] = 80'h0010ffabffabffabffab;
mem[5061] = 80'h0010ffabffabffabffab;
mem[5062] = 80'h0010ffabffabffabffab;
mem[5063] = 80'h0010ffabffabffabffab;
mem[5064] = 80'h0010ffabffabffabffab;
mem[5065] = 80'h0010ffabffabffabffab;
mem[5066] = 80'h0010ffabffabffabffab;
mem[5067] = 80'h0010ffabffabffabffab;
mem[5068] = 80'h0010ffabffabffabffab;
mem[5069] = 80'h0010ffabffabffabffab;
mem[5070] = 80'h0010ffabffabffabffab;
mem[5071] = 80'h0010ffabffabffabffab;
mem[5072] = 80'h0010ffabffabffabffab;
mem[5073] = 80'h0010ffabffabffabffab;
mem[5074] = 80'h0010ffabffabffabffab;
mem[5075] = 80'h0010ffabffabffabffab;
mem[5076] = 80'h0010ffabffabffabffab;
mem[5077] = 80'h0010ffabffabffabffab;
mem[5078] = 80'h0010ffabffabffabffab;
mem[5079] = 80'h0010ffabffabffabffab;
mem[5080] = 80'h0010ffabffabffabffab;
mem[5081] = 80'h0010ffabffabffabffab;
mem[5082] = 80'h0010ffabffabffabffab;
mem[5083] = 80'h0010ffabffabffabffab;
mem[5084] = 80'h0010ffabffabffabffab;
mem[5085] = 80'h0010ffabffabffabffab;
mem[5086] = 80'h0010ffabffabffabffab;
mem[5087] = 80'h0010ffabffabffabffab;
mem[5088] = 80'h0010ffabffabffabffab;
mem[5089] = 80'h0010ffabffabffabffab;
mem[5090] = 80'h0010ffabffabffabffab;
mem[5091] = 80'h0010ffabffabffabffab;
mem[5092] = 80'h0010ffabffabffabffab;
mem[5093] = 80'h0010ffabffabffabffab;
mem[5094] = 80'h0010ffabffabffabffab;
mem[5095] = 80'h0010ffabffabffabffab;
mem[5096] = 80'h0010ffabffabffabffab;
mem[5097] = 80'h0010ffabffabffabffab;
mem[5098] = 80'h0010ffabffabffabffab;
mem[5099] = 80'h0010ffabffabffabffab;
mem[5100] = 80'h0010ffabffabffabffab;
mem[5101] = 80'h0010ffabffabffabffab;
mem[5102] = 80'h0010ffabffabffabffab;
mem[5103] = 80'h0010ffabffabffabffab;
mem[5104] = 80'h0010ffabffabffabffab;
mem[5105] = 80'h0010ffabffabffabffab;
mem[5106] = 80'h0010ffabffabffabffab;
mem[5107] = 80'h0010ffabffabffabffab;
mem[5108] = 80'h0010ffabffabffabffab;
mem[5109] = 80'h0010ffabffabffabffab;
mem[5110] = 80'h0010ffabffabffabffab;
mem[5111] = 80'h0010ffabffabffabffab;
mem[5112] = 80'h0010ffabffabffabffab;
mem[5113] = 80'h0010ffabffabffabffab;
mem[5114] = 80'h0010ffabffabffabffab;
mem[5115] = 80'h0010ffabffabffabffab;
mem[5116] = 80'h0010ffabffabffabffab;
mem[5117] = 80'h0010ffabffabffabffab;
mem[5118] = 80'h0010ffabffabffabffab;
mem[5119] = 80'h0010ffabffabffabffab;
mem[5120] = 80'h0010ffabffabffabffab;
mem[5121] = 80'h0010ffabffabffabffab;
mem[5122] = 80'h0010ffabffabffabffab;
mem[5123] = 80'h0010ffabffabffabffab;
mem[5124] = 80'h0010ffabffabffabffab;
mem[5125] = 80'h0010ffabffabffabffab;
mem[5126] = 80'h0010ffabffabffabffab;
mem[5127] = 80'h0010ffabffabffabffab;
mem[5128] = 80'h0010ffabffabffabffab;
mem[5129] = 80'h0010ffabffabffabffab;
mem[5130] = 80'h0010ffabffabffabffab;
mem[5131] = 80'h0010ffabffabffabffab;
mem[5132] = 80'h0010ffabffabff361e71;
mem[5133] = 80'h0010aff27d29cd0afdd0;
mem[5134] = 80'h001091875471dd9418d3;
mem[5135] = 80'h01150d7b4ab987000000;
mem[5136] = 80'h10100000010000010010;
mem[5137] = 80'h00109400000208004500;
mem[5138] = 80'h0010015c89ca0000fffd;
mem[5139] = 80'h0010ae81c0550102c000;
mem[5140] = 80'h00100001ffabffabffab;
mem[5141] = 80'h0010ffabffabffabffab;
mem[5142] = 80'h0010ffabffabffabffab;
mem[5143] = 80'h0010ffabffabffabffab;
mem[5144] = 80'h0010ffabffabffabffab;
mem[5145] = 80'h0010ffabffabffabffab;
mem[5146] = 80'h0010ffabffabffabffab;
mem[5147] = 80'h0010ffabffabffabffab;
mem[5148] = 80'h0010ffabffabffabffab;
mem[5149] = 80'h0010ffabffabffabffab;
mem[5150] = 80'h0010ffabffabffabffab;
mem[5151] = 80'h0010ffabffabffabffab;
mem[5152] = 80'h0010ffabffabffabffab;
mem[5153] = 80'h0010ffabffabffabffab;
mem[5154] = 80'h0010ffabffabffabffab;
mem[5155] = 80'h0010ffabffabffabffab;
mem[5156] = 80'h0010ffabffabffabffab;
mem[5157] = 80'h0010ffabffabffabffab;
mem[5158] = 80'h0010ffabffabffabffab;
mem[5159] = 80'h0010ffabffabffabffab;
mem[5160] = 80'h0010ffabffabffabffab;
mem[5161] = 80'h0010ffabffabffabffab;
mem[5162] = 80'h0010ffabffabffabffab;
mem[5163] = 80'h0010ffabffabffabffab;
mem[5164] = 80'h0010ffabffabffabffab;
mem[5165] = 80'h0010ffabffabffabffab;
mem[5166] = 80'h0010ffabffabffabffab;
mem[5167] = 80'h0010ffabffabffabffab;
mem[5168] = 80'h0010ffabffabffabffab;
mem[5169] = 80'h0010ffabffabffabffab;
mem[5170] = 80'h0010ffabffabffabffab;
mem[5171] = 80'h0010ffabffabffabffab;
mem[5172] = 80'h0010ffabffabffabffab;
mem[5173] = 80'h0010ffabffabffabffab;
mem[5174] = 80'h0010ffabffabffabffab;
mem[5175] = 80'h0010ffabffabffabffab;
mem[5176] = 80'h0010ffabffabffabffab;
mem[5177] = 80'h0010ffabffabffabffab;
mem[5178] = 80'h0010ffabffabffab358c;
mem[5179] = 80'h001013da9af76e0d568a;
mem[5180] = 80'h001058a79925b82f8d9b;
mem[5181] = 80'h01161f7258a1b0770000;
mem[5182] = 80'h10100000010000010010;
mem[5183] = 80'h00109400000208004500;
mem[5184] = 80'h001000c589cb0000fffd;
mem[5185] = 80'h0010af17c0550102c000;
mem[5186] = 80'h00100001ffabffabffab;
mem[5187] = 80'h0010ffabffabffabffab;
mem[5188] = 80'h0010ffabffabffabffab;
mem[5189] = 80'h0010ffabffabffabffab;
mem[5190] = 80'h0010ffabffabffabffab;
mem[5191] = 80'h0010ffabffabffabffab;
mem[5192] = 80'h0010ffabffabffabffab;
mem[5193] = 80'h0010ffabffabffabffab;
mem[5194] = 80'h0010ffabffabffabffab;
mem[5195] = 80'h0010ffabffabffabffab;
mem[5196] = 80'h0010ffabffabffabffab;
mem[5197] = 80'h0010ffabffabffabffab;
mem[5198] = 80'h0010ffabffabffabffab;
mem[5199] = 80'h0010ffabffabffabffab;
mem[5200] = 80'h0010ffabffabffabffab;
mem[5201] = 80'h0010ffabffabffabffab;
mem[5202] = 80'h0010ffabffabffabffab;
mem[5203] = 80'h0010ffabffabffabffab;
mem[5204] = 80'h0010ffabffabffabffab;
mem[5205] = 80'h0010ffabffabffabff34;
mem[5206] = 80'h0010fdcdf6428eacb29d;
mem[5207] = 80'h001058df4a6cf5417e55;
mem[5208] = 80'h0117088dab6f4e01d100;
mem[5209] = 80'h10100000010000010010;
mem[5210] = 80'h00109400000208004500;
mem[5211] = 80'h0010007889cc0000fffd;
mem[5212] = 80'h0010af63c0550102c000;
mem[5213] = 80'h00100001ffabffabffab;
mem[5214] = 80'h0010ffabffabffabffab;
mem[5215] = 80'h0010ffabffabffabffab;
mem[5216] = 80'h0010ffabffabffabffab;
mem[5217] = 80'h0010ffabffabffabffab;
mem[5218] = 80'h0010ffabffabffabffab;
mem[5219] = 80'h0010ffabffabffabffab;
mem[5220] = 80'h0010ffabffabffabffab;
mem[5221] = 80'h0010ffabffabffabffab;
mem[5222] = 80'h0010ffabffabffabffab;
mem[5223] = 80'h0010ffab33d9091c939a;
mem[5224] = 80'h0010233225b7ce265014;
mem[5225] = 80'h00104a9bccadb102c73a;
mem[5226] = 80'h0112473e000000000000;
mem[5227] = 80'h10100000010000010010;
mem[5228] = 80'h00109400000208004500;
mem[5229] = 80'h0010005389cd0000fffd;
mem[5230] = 80'h0010af87c0550102c000;
mem[5231] = 80'h00100001ffabffabffab;
mem[5232] = 80'h0010ffabffabffabffab;
mem[5233] = 80'h0010ffabffabffabffab;
mem[5234] = 80'h0010ffabffabffabffab;
mem[5235] = 80'h0010ffabffabffabffab;
mem[5236] = 80'h0010ffabffabff32a8d7;
mem[5237] = 80'h0010304be3e18dee6549;
mem[5238] = 80'h0010cba5c7f8ca9c5855;
mem[5239] = 80'h01159961f14d22000000;
mem[5240] = 80'h10100000010000010010;
mem[5241] = 80'h00109400000208004500;
mem[5242] = 80'h0010031889ce0000fffd;
mem[5243] = 80'h0010acc1c0550102c000;
mem[5244] = 80'h00100001ffabffabffab;
mem[5245] = 80'h0010ffabffabffabffab;
mem[5246] = 80'h0010ffabffabffabffab;
mem[5247] = 80'h0010ffabffabffabffab;
mem[5248] = 80'h0010ffabffabffabffab;
mem[5249] = 80'h0010ffabffabffabffab;
mem[5250] = 80'h0010ffabffabffabffab;
mem[5251] = 80'h0010ffabffabffabffab;
mem[5252] = 80'h0010ffabffabffabffab;
mem[5253] = 80'h0010ffabffabffabffab;
mem[5254] = 80'h0010ffabffabffabffab;
mem[5255] = 80'h0010ffabffabffabffab;
mem[5256] = 80'h0010ffabffabffabffab;
mem[5257] = 80'h0010ffabffabffabffab;
mem[5258] = 80'h0010ffabffabffabffab;
mem[5259] = 80'h0010ffabffabffabffab;
mem[5260] = 80'h0010ffabffabffabffab;
mem[5261] = 80'h0010ffabffabffabffab;
mem[5262] = 80'h0010ffabffabffabffab;
mem[5263] = 80'h0010ffabffabffabffab;
mem[5264] = 80'h0010ffabffabffabffab;
mem[5265] = 80'h0010ffabffabffabffab;
mem[5266] = 80'h0010ffabffabffabffab;
mem[5267] = 80'h0010ffabffabffabffab;
mem[5268] = 80'h0010ffabffabffabffab;
mem[5269] = 80'h0010ffabffabffabffab;
mem[5270] = 80'h0010ffabffabffabffab;
mem[5271] = 80'h0010ffabffabffabffab;
mem[5272] = 80'h0010ffabffabffabffab;
mem[5273] = 80'h0010ffabffabffabffab;
mem[5274] = 80'h0010ffabffabffabffab;
mem[5275] = 80'h0010ffabffabffabffab;
mem[5276] = 80'h0010ffabffabffabffab;
mem[5277] = 80'h0010ffabffabffabffab;
mem[5278] = 80'h0010ffabffabffabffab;
mem[5279] = 80'h0010ffabffabffabffab;
mem[5280] = 80'h0010ffabffabffabffab;
mem[5281] = 80'h0010ffabffabffabffab;
mem[5282] = 80'h0010ffabffabffabffab;
mem[5283] = 80'h0010ffabffabffabffab;
mem[5284] = 80'h0010ffabffabffabffab;
mem[5285] = 80'h0010ffabffabffabffab;
mem[5286] = 80'h0010ffabffabffabffab;
mem[5287] = 80'h0010ffabffabffabffab;
mem[5288] = 80'h0010ffabffabffabffab;
mem[5289] = 80'h0010ffabffabffabffab;
mem[5290] = 80'h0010ffabffabffabffab;
mem[5291] = 80'h0010ffabffabffabffab;
mem[5292] = 80'h0010ffabffabffabffab;
mem[5293] = 80'h0010ffabffabffabffab;
mem[5294] = 80'h0010ffabffabffabffab;
mem[5295] = 80'h0010ffabffabffabffab;
mem[5296] = 80'h0010ffabffabffabffab;
mem[5297] = 80'h0010ffabffabffabffab;
mem[5298] = 80'h0010ffabffabffabffab;
mem[5299] = 80'h0010ffabffabffabffab;
mem[5300] = 80'h0010ffabffabffabffab;
mem[5301] = 80'h0010ffabffabffabffab;
mem[5302] = 80'h0010ffabffabffabffab;
mem[5303] = 80'h0010ffabffabffabffab;
mem[5304] = 80'h0010ffabffabffabffab;
mem[5305] = 80'h0010ffabffabffabffab;
mem[5306] = 80'h0010ffabffabffabffab;
mem[5307] = 80'h0010ffabffabffabffab;
mem[5308] = 80'h0010ffabffabffabffab;
mem[5309] = 80'h0010ffabffabffabffab;
mem[5310] = 80'h0010ffabffabffabffab;
mem[5311] = 80'h0010ffabffabffabffab;
mem[5312] = 80'h0010ffabffabffabffab;
mem[5313] = 80'h0010ffabffabffabffab;
mem[5314] = 80'h0010ffabffabffabffab;
mem[5315] = 80'h0010ffabffabffabffab;
mem[5316] = 80'h0010ffabffabffabffab;
mem[5317] = 80'h0010ffabffabffabffab;
mem[5318] = 80'h0010ffabffabffabffab;
mem[5319] = 80'h0010ffabffabffabffab;
mem[5320] = 80'h0010ffabffabffabffab;
mem[5321] = 80'h0010ffabffabffabffab;
mem[5322] = 80'h0010ffabffabffabffab;
mem[5323] = 80'h0010ffabffabffabffab;
mem[5324] = 80'h0010ffabffabffabffab;
mem[5325] = 80'h0010ffabffabffabffab;
mem[5326] = 80'h0010ffabffabffabffab;
mem[5327] = 80'h0010ffabffabffabffab;
mem[5328] = 80'h0010ffabffabffabffab;
mem[5329] = 80'h0010ffabffabffabffab;
mem[5330] = 80'h0010ffabffabffabffab;
mem[5331] = 80'h0010ffabffabffabffab;
mem[5332] = 80'h0010ffabffabffabffab;
mem[5333] = 80'h0010ffabffabffabffab;
mem[5334] = 80'h0010ffabffabffabffab;
mem[5335] = 80'h0010ffabffabffabffab;
mem[5336] = 80'h0010ffabffabffabffab;
mem[5337] = 80'h0010ffabffabffabffab;
mem[5338] = 80'h0010ffab313ab5452369;
mem[5339] = 80'h0010a64db212c1fdbbb7;
mem[5340] = 80'h00102e38a1a650226991;
mem[5341] = 80'h01129bfe000000000000;
mem[5342] = 80'h10100000010000010010;
mem[5343] = 80'h00109400000208004500;
mem[5344] = 80'h0010047a89cf0000fffd;
mem[5345] = 80'h0010ab5ec0550102c000;
mem[5346] = 80'h00100001ffabffabffab;
mem[5347] = 80'h0010ffabffabffabffab;
mem[5348] = 80'h0010ffabffabffabffab;
mem[5349] = 80'h0010ffabffabffabffab;
mem[5350] = 80'h0010ffabffabffabffab;
mem[5351] = 80'h0010ffabffabffabffab;
mem[5352] = 80'h0010ffabffabffabffab;
mem[5353] = 80'h0010ffabffabffabffab;
mem[5354] = 80'h0010ffabffabffabffab;
mem[5355] = 80'h0010ffabffabffabffab;
mem[5356] = 80'h0010ffabffabffabffab;
mem[5357] = 80'h0010ffabffabffabffab;
mem[5358] = 80'h0010ffabffabffabffab;
mem[5359] = 80'h0010ffabffabffabffab;
mem[5360] = 80'h0010ffabffabffabffab;
mem[5361] = 80'h0010ffabffabffabffab;
mem[5362] = 80'h0010ffabffabffabffab;
mem[5363] = 80'h0010ffabffabffabffab;
mem[5364] = 80'h0010ffabffabffabffab;
mem[5365] = 80'h0010ffabffabffabffab;
mem[5366] = 80'h0010ffabffabffabffab;
mem[5367] = 80'h0010ffabffabffabffab;
mem[5368] = 80'h0010ffabffabffabffab;
mem[5369] = 80'h0010ffabffabffabffab;
mem[5370] = 80'h0010ffabffabffabffab;
mem[5371] = 80'h0010ffabffabffabffab;
mem[5372] = 80'h0010ffabffabffabffab;
mem[5373] = 80'h0010ffabffabffabffab;
mem[5374] = 80'h0010ffabffabffabffab;
mem[5375] = 80'h0010ffabffabffabffab;
mem[5376] = 80'h0010ffabffabffabffab;
mem[5377] = 80'h0010ffabffabffabffab;
mem[5378] = 80'h0010ffabffabffabffab;
mem[5379] = 80'h0010ffabffabffabffab;
mem[5380] = 80'h0010ffabffabffabffab;
mem[5381] = 80'h0010ffabffabffabffab;
mem[5382] = 80'h0010ffabffabffabffab;
mem[5383] = 80'h0010ffabffabffabffab;
mem[5384] = 80'h0010ffabffabffabffab;
mem[5385] = 80'h0010ffabffabffabffab;
mem[5386] = 80'h0010ffabffabffabffab;
mem[5387] = 80'h0010ffabffabffabffab;
mem[5388] = 80'h0010ffabffabffabffab;
mem[5389] = 80'h0010ffabffabffabffab;
mem[5390] = 80'h0010ffabffabffabffab;
mem[5391] = 80'h0010ffabffabffabffab;
mem[5392] = 80'h0010ffabffabffabffab;
mem[5393] = 80'h0010ffabffabffabffab;
mem[5394] = 80'h0010ffabffabffabffab;
mem[5395] = 80'h0010ffabffabffabffab;
mem[5396] = 80'h0010ffabffabffabffab;
mem[5397] = 80'h0010ffabffabffabffab;
mem[5398] = 80'h0010ffabffabffabffab;
mem[5399] = 80'h0010ffabffabffabffab;
mem[5400] = 80'h0010ffabffabffabffab;
mem[5401] = 80'h0010ffabffabffabffab;
mem[5402] = 80'h0010ffabffabffabffab;
mem[5403] = 80'h0010ffabffabffabffab;
mem[5404] = 80'h0010ffabffabffabffab;
mem[5405] = 80'h0010ffabffabffabffab;
mem[5406] = 80'h0010ffabffabffabffab;
mem[5407] = 80'h0010ffabffabffabffab;
mem[5408] = 80'h0010ffabffabffabffab;
mem[5409] = 80'h0010ffabffabffabffab;
mem[5410] = 80'h0010ffabffabffabffab;
mem[5411] = 80'h0010ffabffabffabffab;
mem[5412] = 80'h0010ffabffabffabffab;
mem[5413] = 80'h0010ffabffabffabffab;
mem[5414] = 80'h0010ffabffabffabffab;
mem[5415] = 80'h0010ffabffabffabffab;
mem[5416] = 80'h0010ffabffabffabffab;
mem[5417] = 80'h0010ffabffabffabffab;
mem[5418] = 80'h0010ffabffabffabffab;
mem[5419] = 80'h0010ffabffabffabffab;
mem[5420] = 80'h0010ffabffabffabffab;
mem[5421] = 80'h0010ffabffabffabffab;
mem[5422] = 80'h0010ffabffabffabffab;
mem[5423] = 80'h0010ffabffabffabffab;
mem[5424] = 80'h0010ffabffabffabffab;
mem[5425] = 80'h0010ffabffabffabffab;
mem[5426] = 80'h0010ffabffabffabffab;
mem[5427] = 80'h0010ffabffabffabffab;
mem[5428] = 80'h0010ffabffabffabffab;
mem[5429] = 80'h0010ffabffabffabffab;
mem[5430] = 80'h0010ffabffabffabffab;
mem[5431] = 80'h0010ffabffabffabffab;
mem[5432] = 80'h0010ffabffabffabffab;
mem[5433] = 80'h0010ffabffabffabffab;
mem[5434] = 80'h0010ffabffabffabffab;
mem[5435] = 80'h0010ffabffabffabffab;
mem[5436] = 80'h0010ffabffabffabffab;
mem[5437] = 80'h0010ffabffabffabffab;
mem[5438] = 80'h0010ffabffabffabffab;
mem[5439] = 80'h0010ffabffabffabffab;
mem[5440] = 80'h0010ffabffabffabffab;
mem[5441] = 80'h0010ffabffabffabffab;
mem[5442] = 80'h0010ffabffabffabffab;
mem[5443] = 80'h0010ffabffabffabffab;
mem[5444] = 80'h0010ffabffabffabffab;
mem[5445] = 80'h0010ffabffabffabffab;
mem[5446] = 80'h0010ffabffabffabffab;
mem[5447] = 80'h0010ffabffabffabffab;
mem[5448] = 80'h0010ffabffabffabffab;
mem[5449] = 80'h0010ffabffabffabffab;
mem[5450] = 80'h0010ffabffabffabffab;
mem[5451] = 80'h0010ffabffabffabffab;
mem[5452] = 80'h0010ffabffabffabffab;
mem[5453] = 80'h0010ffabffabffabffab;
mem[5454] = 80'h0010ffabffabffabffab;
mem[5455] = 80'h0010ffabffabffabffab;
mem[5456] = 80'h0010ffabffabffabffab;
mem[5457] = 80'h0010ffabffabffabffab;
mem[5458] = 80'h0010ffabffabffabffab;
mem[5459] = 80'h0010ffabffabffabffab;
mem[5460] = 80'h0010ffabffabffabffab;
mem[5461] = 80'h0010ffabffabffabffab;
mem[5462] = 80'h0010ffabffabffabffab;
mem[5463] = 80'h0010ffabffabffabffab;
mem[5464] = 80'h0010ffabffabffabffab;
mem[5465] = 80'h0010ffabffabffabffab;
mem[5466] = 80'h0010ffabffabffabffab;
mem[5467] = 80'h0010ffabffabffabffab;
mem[5468] = 80'h0010ffabffabffabffab;
mem[5469] = 80'h0010ffabffabffabffab;
mem[5470] = 80'h0010ffabffabffabffab;
mem[5471] = 80'h0010ffabffabffabffab;
mem[5472] = 80'h0010ffabffabffabffab;
mem[5473] = 80'h0010ffabffabffabffab;
mem[5474] = 80'h0010ffabffabffabffab;
mem[5475] = 80'h0010ffabffabffabffab;
mem[5476] = 80'h0010ffabffabffabffab;
mem[5477] = 80'h0010ffabffabffabffab;
mem[5478] = 80'h0010ffabffabffabffab;
mem[5479] = 80'h0010ffabffabffabffab;
mem[5480] = 80'h0010ffabffabffabffab;
mem[5481] = 80'h0010ffabffabffabffab;
mem[5482] = 80'h0010ffabffabffabffab;
mem[5483] = 80'h0010ffabffabffabffab;
mem[5484] = 80'h0010ffabffab304b6b69;
mem[5485] = 80'h0010fb1064f279c04610;
mem[5486] = 80'h00104e664169fc48b85e;
mem[5487] = 80'h011441bc72fd00000000;
mem[5488] = 80'h00000000000000000000;
mem[5489] = 80'h00000000000000000000;
mem[5490] = 80'h00000000000000000000;
mem[5491] = 80'h00000000000000000000;
mem[5492] = 80'h00000000000000000000;
mem[5493] = 80'h00000000000000000000;
mem[5494] = 80'h00000000000000000000;
mem[5495] = 80'h00000000000000000000;
mem[5496] = 80'h00000000000000000000;
mem[5497] = 80'h00000000000000000000;
mem[5498] = 80'h00000000000000000000;
mem[5499] = 80'h00000000000000000000;
mem[5500] = 80'h00000000000000000000;
mem[5501] = 80'h00000000000000000000;
mem[5502] = 80'h00000000000000000000;
mem[5503] = 80'h00000000000000000000;
mem[5504] = 80'h00000000000000000000;
mem[5505] = 80'h00000000000000000000;
mem[5506] = 80'h00000000000000000000;
mem[5507] = 80'h00000000000000000000;
mem[5508] = 80'h00000000000000000000;
mem[5509] = 80'h00000000000000000000;
mem[5510] = 80'h00000000000000000000;
mem[5511] = 80'h00000000000000000000;
mem[5512] = 80'h00000000000000000000;
mem[5513] = 80'h10100000010000010010;
mem[5514] = 80'h00109400000208004500;
mem[5515] = 80'h0010052b89d00000fffd;
mem[5516] = 80'h0010aaacc0550102c000;
mem[5517] = 80'h00100001ffabffabffab;
mem[5518] = 80'h0010ffabffabffabffab;
mem[5519] = 80'h0010ffabffabffabffab;
mem[5520] = 80'h0010ffabffabffabffab;
mem[5521] = 80'h0010ffabffabffabffab;
mem[5522] = 80'h0010ffabffabffabffab;
mem[5523] = 80'h0010ffabffabffabffab;
mem[5524] = 80'h0010ffabffabffabffab;
mem[5525] = 80'h0010ffabffabffabffab;
mem[5526] = 80'h0010ffabffabffabffab;
mem[5527] = 80'h0010ffabffabffabffab;
mem[5528] = 80'h0010ffabffabffabffab;
mem[5529] = 80'h0010ffabffabffabffab;
mem[5530] = 80'h0010ffabffabffabffab;
mem[5531] = 80'h0010ffabffabffabffab;
mem[5532] = 80'h0010ffabffabffabffab;
mem[5533] = 80'h0010ffabffabffabffab;
mem[5534] = 80'h0010ffabffabffabffab;
mem[5535] = 80'h0010ffabffabffabffab;
mem[5536] = 80'h0010ffabffabffabffab;
mem[5537] = 80'h0010ffabffabffabffab;
mem[5538] = 80'h0010ffabffabffabffab;
mem[5539] = 80'h0010ffabffabffabffab;
mem[5540] = 80'h0010ffabffabffabffab;
mem[5541] = 80'h0010ffabffabffabffab;
mem[5542] = 80'h0010ffabffabffabffab;
mem[5543] = 80'h0010ffabffabffabffab;
mem[5544] = 80'h0010ffabffabffabffab;
mem[5545] = 80'h0010ffabffabffabffab;
mem[5546] = 80'h0010ffabffabffabffab;
mem[5547] = 80'h0010ffabffabffabffab;
mem[5548] = 80'h0010ffabffabffabffab;
mem[5549] = 80'h0010ffabffabffabffab;
mem[5550] = 80'h0010ffabffabffabffab;
mem[5551] = 80'h0010ffabffabffabffab;
mem[5552] = 80'h0010ffabffabffabffab;
mem[5553] = 80'h0010ffabffabffabffab;
mem[5554] = 80'h0010ffabffabffabffab;
mem[5555] = 80'h0010ffabffabffabffab;
mem[5556] = 80'h0010ffabffabffabffab;
mem[5557] = 80'h0010ffabffabffabffab;
mem[5558] = 80'h0010ffabffabffabffab;
mem[5559] = 80'h0010ffabffabffabffab;
mem[5560] = 80'h0010ffabffabffabffab;
mem[5561] = 80'h0010ffabffabffabffab;
mem[5562] = 80'h0010ffabffabffabffab;
mem[5563] = 80'h0010ffabffabffabffab;
mem[5564] = 80'h0010ffabffabffabffab;
mem[5565] = 80'h0010ffabffabffabffab;
mem[5566] = 80'h0010ffabffabffabffab;
mem[5567] = 80'h0010ffabffabffabffab;
mem[5568] = 80'h0010ffabffabffabffab;
mem[5569] = 80'h0010ffabffabffabffab;
mem[5570] = 80'h0010ffabffabffabffab;
mem[5571] = 80'h0010ffabffabffabffab;
mem[5572] = 80'h0010ffabffabffabffab;
mem[5573] = 80'h0010ffabffabffabffab;
mem[5574] = 80'h0010ffabffabffabffab;
mem[5575] = 80'h0010ffabffabffabffab;
mem[5576] = 80'h0010ffabffabffabffab;
mem[5577] = 80'h0010ffabffabffabffab;
mem[5578] = 80'h0010ffabffabffabffab;
mem[5579] = 80'h0010ffabffabffabffab;
mem[5580] = 80'h0010ffabffabffabffab;
mem[5581] = 80'h0010ffabffabffabffab;
mem[5582] = 80'h0010ffabffabffabffab;
mem[5583] = 80'h0010ffabffabffabffab;
mem[5584] = 80'h0010ffabffabffabffab;
mem[5585] = 80'h0010ffabffabffabffab;
mem[5586] = 80'h0010ffabffabffabffab;
mem[5587] = 80'h0010ffabffabffabffab;
mem[5588] = 80'h0010ffabffabffabffab;
mem[5589] = 80'h0010ffabffabffabffab;
mem[5590] = 80'h0010ffabffabffabffab;
mem[5591] = 80'h0010ffabffabffabffab;
mem[5592] = 80'h0010ffabffabffabffab;
mem[5593] = 80'h0010ffabffabffabffab;
mem[5594] = 80'h0010ffabffabffabffab;
mem[5595] = 80'h0010ffabffabffabffab;
mem[5596] = 80'h0010ffabffabffabffab;
mem[5597] = 80'h0010ffabffabffabffab;
mem[5598] = 80'h0010ffabffabffabffab;
mem[5599] = 80'h0010ffabffabffabffab;
mem[5600] = 80'h0010ffabffabffabffab;
mem[5601] = 80'h0010ffabffabffabffab;
mem[5602] = 80'h0010ffabffabffabffab;
mem[5603] = 80'h0010ffabffabffabffab;
mem[5604] = 80'h0010ffabffabffabffab;
mem[5605] = 80'h0010ffabffabffabffab;
mem[5606] = 80'h0010ffabffabffabffab;
mem[5607] = 80'h0010ffabffabffabffab;
mem[5608] = 80'h0010ffabffabffabffab;
mem[5609] = 80'h0010ffabffabffabffab;
mem[5610] = 80'h0010ffabffabffabffab;
mem[5611] = 80'h0010ffabffabffabffab;
mem[5612] = 80'h0010ffabffabffabffab;
mem[5613] = 80'h0010ffabffabffabffab;
mem[5614] = 80'h0010ffabffabffabffab;
mem[5615] = 80'h0010ffabffabffabffab;
mem[5616] = 80'h0010ffabffabffabffab;
mem[5617] = 80'h0010ffabffabffabffab;
mem[5618] = 80'h0010ffabffabffabffab;
mem[5619] = 80'h0010ffabffabffabffab;
mem[5620] = 80'h0010ffabffabffabffab;
mem[5621] = 80'h0010ffabffabffabffab;
mem[5622] = 80'h0010ffabffabffabffab;
mem[5623] = 80'h0010ffabffabffabffab;
mem[5624] = 80'h0010ffabffabffabffab;
mem[5625] = 80'h0010ffabffabffabffab;
mem[5626] = 80'h0010ffabffabffabffab;
mem[5627] = 80'h0010ffabffabffabffab;
mem[5628] = 80'h0010ffabffabffabffab;
mem[5629] = 80'h0010ffabffabffabffab;
mem[5630] = 80'h0010ffabffabffabffab;
mem[5631] = 80'h0010ffabffabffabffab;
mem[5632] = 80'h0010ffabffabffabffab;
mem[5633] = 80'h0010ffabffabffabffab;
mem[5634] = 80'h0010ffabffabffabffab;
mem[5635] = 80'h0010ffabffabffabffab;
mem[5636] = 80'h0010ffabffabffabffab;
mem[5637] = 80'h0010ffabffabffabffab;
mem[5638] = 80'h0010ffabffabffabffab;
mem[5639] = 80'h0010ffabffabffabffab;
mem[5640] = 80'h0010ffabffabffabffab;
mem[5641] = 80'h0010ffabffabffabffab;
mem[5642] = 80'h0010ffabffabffabffab;
mem[5643] = 80'h0010ffabffabffabffab;
mem[5644] = 80'h0010ffabffabffabffab;
mem[5645] = 80'h0010ffabffabffabffab;
mem[5646] = 80'h0010ffabffabffabffab;
mem[5647] = 80'h0010ffabffabffabffab;
mem[5648] = 80'h0010ffabffabffabffab;
mem[5649] = 80'h0010ffabffabffabffab;
mem[5650] = 80'h0010ffabffabffabffab;
mem[5651] = 80'h0010ffabffabffabffab;
mem[5652] = 80'h0010ffabffabffabffab;
mem[5653] = 80'h0010ffabffabffabffab;
mem[5654] = 80'h0010ffabffabffabffab;
mem[5655] = 80'h0010ffabffabffabffab;
mem[5656] = 80'h0010ffabffabffabffab;
mem[5657] = 80'h0010ffabffabffabffab;
mem[5658] = 80'h0010ffabffabffabffab;
mem[5659] = 80'h0010ffabffabffabffab;
mem[5660] = 80'h0010ffabffabffabffab;
mem[5661] = 80'h0010ffabffabffabffab;
mem[5662] = 80'h0010ffabffabffabffab;
mem[5663] = 80'h0010ffabffabffabffab;
mem[5664] = 80'h0010ffabffabffabffab;
mem[5665] = 80'h0010ffabffabffabffab;
mem[5666] = 80'h0010ffabffabffabffab;
mem[5667] = 80'h0010ffabffabffabffab;
mem[5668] = 80'h0010ffabffabffabffab;
mem[5669] = 80'h0010ffabffabffabffab;
mem[5670] = 80'h0010ffabffabffabffab;
mem[5671] = 80'h0010ffabffabffabffab;
mem[5672] = 80'h0010ffabffabffabffab;
mem[5673] = 80'h0010ffabffabffabffab;
mem[5674] = 80'h0010ffabffabffabffab;
mem[5675] = 80'h0010ffabffabffabffab;
mem[5676] = 80'h0010ffabffabffabffab;
mem[5677] = 80'h0010ffabffabff2f4a1a;
mem[5678] = 80'h0010b7d7c81d30c60b8b;
mem[5679] = 80'h001096a38c160cd110e4;
mem[5680] = 80'h0115b95a12d171000000;
mem[5681] = 80'h00000000000000000000;
mem[5682] = 80'h00000000000000000000;
mem[5683] = 80'h00000000000000000000;
mem[5684] = 80'h00000000000000000000;
mem[5685] = 80'h00000000000000000000;
mem[5686] = 80'h00000000000000000000;
mem[5687] = 80'h00000000000000000000;
mem[5688] = 80'h00000000000000000000;
mem[5689] = 80'h00000000000000000000;
mem[5690] = 80'h00000000000000000000;
mem[5691] = 80'h00000000000000000000;
mem[5692] = 80'h00000000000000000000;
mem[5693] = 80'h00000000000000000000;
mem[5694] = 80'h00000000000000000000;
mem[5695] = 80'h10100000010000010010;
mem[5696] = 80'h00109400000208004500;
mem[5697] = 80'h0010058389d10000fffd;
mem[5698] = 80'h0010aa53c0550102c000;
mem[5699] = 80'h00100001ffabffabffab;
mem[5700] = 80'h0010ffabffabffabffab;
mem[5701] = 80'h0010ffabffabffabffab;
mem[5702] = 80'h0010ffabffabffabffab;
mem[5703] = 80'h0010ffabffabffabffab;
mem[5704] = 80'h0010ffabffabffabffab;
mem[5705] = 80'h0010ffabffabffabffab;
mem[5706] = 80'h0010ffabffabffabffab;
mem[5707] = 80'h0010ffabffabffabffab;
mem[5708] = 80'h0010ffabffabffabffab;
mem[5709] = 80'h0010ffabffabffabffab;
mem[5710] = 80'h0010ffabffabffabffab;
mem[5711] = 80'h0010ffabffabffabffab;
mem[5712] = 80'h0010ffabffabffabffab;
mem[5713] = 80'h0010ffabffabffabffab;
mem[5714] = 80'h0010ffabffabffabffab;
mem[5715] = 80'h0010ffabffabffabffab;
mem[5716] = 80'h0010ffabffabffabffab;
mem[5717] = 80'h0010ffabffabffabffab;
mem[5718] = 80'h0010ffabffabffabffab;
mem[5719] = 80'h0010ffabffabffabffab;
mem[5720] = 80'h0010ffabffabffabffab;
mem[5721] = 80'h0010ffabffabffabffab;
mem[5722] = 80'h0010ffabffabffabffab;
mem[5723] = 80'h0010ffabffabffabffab;
mem[5724] = 80'h0010ffabffabffabffab;
mem[5725] = 80'h0010ffabffabffabffab;
mem[5726] = 80'h0010ffabffabffabffab;
mem[5727] = 80'h0010ffabffabffabffab;
mem[5728] = 80'h0010ffabffabffabffab;
mem[5729] = 80'h0010ffabffabffabffab;
mem[5730] = 80'h0010ffabffabffabffab;
mem[5731] = 80'h0010ffabffabffabffab;
mem[5732] = 80'h0010ffabffabffabffab;
mem[5733] = 80'h0010ffabffabffabffab;
mem[5734] = 80'h0010ffabffabffabffab;
mem[5735] = 80'h0010ffabffabffabffab;
mem[5736] = 80'h0010ffabffabffabffab;
mem[5737] = 80'h0010ffabffabffabffab;
mem[5738] = 80'h0010ffabffabffabffab;
mem[5739] = 80'h0010ffabffabffabffab;
mem[5740] = 80'h0010ffabffabffabffab;
mem[5741] = 80'h0010ffabffabffabffab;
mem[5742] = 80'h0010ffabffabffabffab;
mem[5743] = 80'h0010ffabffabffabffab;
mem[5744] = 80'h0010ffabffabffabffab;
mem[5745] = 80'h0010ffabffabffabffab;
mem[5746] = 80'h0010ffabffabffabffab;
mem[5747] = 80'h0010ffabffabffabffab;
mem[5748] = 80'h0010ffabffabffabffab;
mem[5749] = 80'h0010ffabffabffabffab;
mem[5750] = 80'h0010ffabffabffabffab;
mem[5751] = 80'h0010ffabffabffabffab;
mem[5752] = 80'h0010ffabffabffabffab;
mem[5753] = 80'h0010ffabffabffabffab;
mem[5754] = 80'h0010ffabffabffabffab;
mem[5755] = 80'h0010ffabffabffabffab;
mem[5756] = 80'h0010ffabffabffabffab;
mem[5757] = 80'h0010ffabffabffabffab;
mem[5758] = 80'h0010ffabffabffabffab;
mem[5759] = 80'h0010ffabffabffabffab;
mem[5760] = 80'h0010ffabffabffabffab;
mem[5761] = 80'h0010ffabffabffabffab;
mem[5762] = 80'h0010ffabffabffabffab;
mem[5763] = 80'h0010ffabffabffabffab;
mem[5764] = 80'h0010ffabffabffabffab;
mem[5765] = 80'h0010ffabffabffabffab;
mem[5766] = 80'h0010ffabffabffabffab;
mem[5767] = 80'h0010ffabffabffabffab;
mem[5768] = 80'h0010ffabffabffabffab;
mem[5769] = 80'h0010ffabffabffabffab;
mem[5770] = 80'h0010ffabffabffabffab;
mem[5771] = 80'h0010ffabffabffabffab;
mem[5772] = 80'h0010ffabffabffabffab;
mem[5773] = 80'h0010ffabffabffabffab;
mem[5774] = 80'h0010ffabffabffabffab;
mem[5775] = 80'h0010ffabffabffabffab;
mem[5776] = 80'h0010ffabffabffabffab;
mem[5777] = 80'h0010ffabffabffabffab;
mem[5778] = 80'h0010ffabffabffabffab;
mem[5779] = 80'h0010ffabffabffabffab;
mem[5780] = 80'h0010ffabffabffabffab;
mem[5781] = 80'h0010ffabffabffabffab;
mem[5782] = 80'h0010ffabffabffabffab;
mem[5783] = 80'h0010ffabffabffabffab;
mem[5784] = 80'h0010ffabffabffabffab;
mem[5785] = 80'h0010ffabffabffabffab;
mem[5786] = 80'h0010ffabffabffabffab;
mem[5787] = 80'h0010ffabffabffabffab;
mem[5788] = 80'h0010ffabffabffabffab;
mem[5789] = 80'h0010ffabffabffabffab;
mem[5790] = 80'h0010ffabffabffabffab;
mem[5791] = 80'h0010ffabffabffabffab;
mem[5792] = 80'h0010ffabffabffabffab;
mem[5793] = 80'h0010ffabffabffabffab;
mem[5794] = 80'h0010ffabffabffabffab;
mem[5795] = 80'h0010ffabffabffabffab;
mem[5796] = 80'h0010ffabffabffabffab;
mem[5797] = 80'h0010ffabffabffabffab;
mem[5798] = 80'h0010ffabffabffabffab;
mem[5799] = 80'h0010ffabffabffabffab;
mem[5800] = 80'h0010ffabffabffabffab;
mem[5801] = 80'h0010ffabffabffabffab;
mem[5802] = 80'h0010ffabffabffabffab;
mem[5803] = 80'h0010ffabffabffabffab;
mem[5804] = 80'h0010ffabffabffabffab;
mem[5805] = 80'h0010ffabffabffabffab;
mem[5806] = 80'h0010ffabffabffabffab;
mem[5807] = 80'h0010ffabffabffabffab;
mem[5808] = 80'h0010ffabffabffabffab;
mem[5809] = 80'h0010ffabffabffabffab;
mem[5810] = 80'h0010ffabffabffabffab;
mem[5811] = 80'h0010ffabffabffabffab;
mem[5812] = 80'h0010ffabffabffabffab;
mem[5813] = 80'h0010ffabffabffabffab;
mem[5814] = 80'h0010ffabffabffabffab;
mem[5815] = 80'h0010ffabffabffabffab;
mem[5816] = 80'h0010ffabffabffabffab;
mem[5817] = 80'h0010ffabffabffabffab;
mem[5818] = 80'h0010ffabffabffabffab;
mem[5819] = 80'h0010ffabffabffabffab;
mem[5820] = 80'h0010ffabffabffabffab;
mem[5821] = 80'h0010ffabffabffabffab;
mem[5822] = 80'h0010ffabffabffabffab;
mem[5823] = 80'h0010ffabffabffabffab;
mem[5824] = 80'h0010ffabffabffabffab;
mem[5825] = 80'h0010ffabffabffabffab;
mem[5826] = 80'h0010ffabffabffabffab;
mem[5827] = 80'h0010ffabffabffabffab;
mem[5828] = 80'h0010ffabffabffabffab;
mem[5829] = 80'h0010ffabffabffabffab;
mem[5830] = 80'h0010ffabffabffabffab;
mem[5831] = 80'h0010ffabffabffabffab;
mem[5832] = 80'h0010ffabffabffabffab;
mem[5833] = 80'h0010ffabffabffabffab;
mem[5834] = 80'h0010ffabffabffabffab;
mem[5835] = 80'h0010ffabffabffabffab;
mem[5836] = 80'h0010ffabffabffabffab;
mem[5837] = 80'h0010ffabffabffabffab;
mem[5838] = 80'h0010ffabffabffabffab;
mem[5839] = 80'h0010ffabffabffabffab;
mem[5840] = 80'h0010ffabffabffabffab;
mem[5841] = 80'h0010ffabffabffabffab;
mem[5842] = 80'h0010ffabffabffabffab;
mem[5843] = 80'h0010ffabffabffabffab;
mem[5844] = 80'h0010ffabffabffabffab;
mem[5845] = 80'h0010ffabffabffabffab;
mem[5846] = 80'h0010ffabffabffabffab;
mem[5847] = 80'h0010ffabffabffabffab;
mem[5848] = 80'h0010ffabffabffabffab;
mem[5849] = 80'h0010ffabffabffabffab;
mem[5850] = 80'h0010ffabffabffabffab;
mem[5851] = 80'h0010ffabffabffabffab;
mem[5852] = 80'h0010ffabffabffabffab;
mem[5853] = 80'h0010ffabffabffabffab;
mem[5854] = 80'h0010ffabffabffabffab;
mem[5855] = 80'h0010ffabffabffabffab;
mem[5856] = 80'h0010ffabffabffabffab;
mem[5857] = 80'h0010ffabffabffabffab;
mem[5858] = 80'h0010ffabffabffabffab;
mem[5859] = 80'h0010ffabffabffabffab;
mem[5860] = 80'h0010ffabffabffabffab;
mem[5861] = 80'h0010ffabffabffabffab;
mem[5862] = 80'h0010ffabffabffabffab;
mem[5863] = 80'h0010ffabffabffabffab;
mem[5864] = 80'h0010ffabffabffabffab;
mem[5865] = 80'h0010ffabffabffabffab;
mem[5866] = 80'h0010ffabffabffabffab;
mem[5867] = 80'h0010ffabffabffabffab;
mem[5868] = 80'h0010ffabffabffabffab;
mem[5869] = 80'h0010ffabffabffabffab;
mem[5870] = 80'h0010ffabffabff2e3bc4;
mem[5871] = 80'h00109b0fb1df8f0dd90c;
mem[5872] = 80'h00107b565e245dad4ddb;
mem[5873] = 80'h01158a53e7b444000000;
mem[5874] = 80'h10100000010000010010;
mem[5875] = 80'h00109400000208004500;
mem[5876] = 80'h001002d989d20000fffd;
mem[5877] = 80'h0010acfcc0550102c000;
mem[5878] = 80'h00100001ffabffabffab;
mem[5879] = 80'h0010ffabffabffabffab;
mem[5880] = 80'h0010ffabffabffabffab;
mem[5881] = 80'h0010ffabffabffabffab;
mem[5882] = 80'h0010ffabffabffabffab;
mem[5883] = 80'h0010ffabffabffabffab;
mem[5884] = 80'h0010ffabffabffabffab;
mem[5885] = 80'h0010ffabffabffabffab;
mem[5886] = 80'h0010ffabffabffabffab;
mem[5887] = 80'h0010ffabffabffabffab;
mem[5888] = 80'h0010ffabffabffabffab;
mem[5889] = 80'h0010ffabffabffabffab;
mem[5890] = 80'h0010ffabffabffabffab;
mem[5891] = 80'h0010ffabffabffabffab;
mem[5892] = 80'h0010ffabffabffabffab;
mem[5893] = 80'h0010ffabffabffabffab;
mem[5894] = 80'h0010ffabffabffabffab;
mem[5895] = 80'h0010ffabffabffabffab;
mem[5896] = 80'h0010ffabffabffabffab;
mem[5897] = 80'h0010ffabffabffabffab;
mem[5898] = 80'h0010ffabffabffabffab;
mem[5899] = 80'h0010ffabffabffabffab;
mem[5900] = 80'h0010ffabffabffabffab;
mem[5901] = 80'h0010ffabffabffabffab;
mem[5902] = 80'h0010ffabffabffabffab;
mem[5903] = 80'h0010ffabffabffabffab;
mem[5904] = 80'h0010ffabffabffabffab;
mem[5905] = 80'h0010ffabffabffabffab;
mem[5906] = 80'h0010ffabffabffabffab;
mem[5907] = 80'h0010ffabffabffabffab;
mem[5908] = 80'h0010ffabffabffabffab;
mem[5909] = 80'h0010ffabffabffabffab;
mem[5910] = 80'h0010ffabffabffabffab;
mem[5911] = 80'h0010ffabffabffabffab;
mem[5912] = 80'h0010ffabffabffabffab;
mem[5913] = 80'h0010ffabffabffabffab;
mem[5914] = 80'h0010ffabffabffabffab;
mem[5915] = 80'h0010ffabffabffabffab;
mem[5916] = 80'h0010ffabffabffabffab;
mem[5917] = 80'h0010ffabffabffabffab;
mem[5918] = 80'h0010ffabffabffabffab;
mem[5919] = 80'h0010ffabffabffabffab;
mem[5920] = 80'h0010ffabffabffabffab;
mem[5921] = 80'h0010ffabffabffabffab;
mem[5922] = 80'h0010ffabffabffabffab;
mem[5923] = 80'h0010ffabffabffabffab;
mem[5924] = 80'h0010ffabffabffabffab;
mem[5925] = 80'h0010ffabffabffabffab;
mem[5926] = 80'h0010ffabffabffabffab;
mem[5927] = 80'h0010ffabffabffabffab;
mem[5928] = 80'h0010ffabffabffabffab;
mem[5929] = 80'h0010ffabffabffabffab;
mem[5930] = 80'h0010ffabffabffabffab;
mem[5931] = 80'h0010ffabffabffabffab;
mem[5932] = 80'h0010ffabffabffabffab;
mem[5933] = 80'h0010ffabffabffabffab;
mem[5934] = 80'h0010ffabffabffabffab;
mem[5935] = 80'h0010ffabffabffabffab;
mem[5936] = 80'h0010ffabffabffabffab;
mem[5937] = 80'h0010ffabffabffabffab;
mem[5938] = 80'h0010ffabffabffabffab;
mem[5939] = 80'h0010ffabffabffabffab;
mem[5940] = 80'h0010ffabffabffabffab;
mem[5941] = 80'h0010ffabffabffabffab;
mem[5942] = 80'h0010ffabffabffabffab;
mem[5943] = 80'h0010ffabffabffabffab;
mem[5944] = 80'h0010ffabffabffabffab;
mem[5945] = 80'h0010ffabffabffabffab;
mem[5946] = 80'h0010ffabffabffabffab;
mem[5947] = 80'h0010ffabffabffabffab;
mem[5948] = 80'h0010ffabffabffabffab;
mem[5949] = 80'h0010ffabffabffabffab;
mem[5950] = 80'h0010ffabffabffabffab;
mem[5951] = 80'h0010ffabffabffabffab;
mem[5952] = 80'h0010ffabffabffabffab;
mem[5953] = 80'h0010ffabffabffabffab;
mem[5954] = 80'h0010ffabffabffabffab;
mem[5955] = 80'h0010ffabffabffabffab;
mem[5956] = 80'h0010ffabffabffabffab;
mem[5957] = 80'h0010ffabffabffabffab;
mem[5958] = 80'h0010ffabffabffabffab;
mem[5959] = 80'h0010ffabffabffabffab;
mem[5960] = 80'h0010ffabffabffabffab;
mem[5961] = 80'h0010ffabffabffabffab;
mem[5962] = 80'h0010ffabffabffabffab;
mem[5963] = 80'h0010ffabffabffabffab;
mem[5964] = 80'h0010ffabff2da9a6ee67;
mem[5965] = 80'h00103b984f51ae844d48;
mem[5966] = 80'h0010285baf85f52c1443;
mem[5967] = 80'h0113924a230000000000;
mem[5968] = 80'h10100000010000010010;
mem[5969] = 80'h00109400000208004500;
mem[5970] = 80'h0010018389d30000fffd;
mem[5971] = 80'h0010ae51c0550102c000;
mem[5972] = 80'h00100001ffabffabffab;
mem[5973] = 80'h0010ffabffabffabffab;
mem[5974] = 80'h0010ffabffabffabffab;
mem[5975] = 80'h0010ffabffabffabffab;
mem[5976] = 80'h0010ffabffabffabffab;
mem[5977] = 80'h0010ffabffabffabffab;
mem[5978] = 80'h0010ffabffabffabffab;
mem[5979] = 80'h0010ffabffabffabffab;
mem[5980] = 80'h0010ffabffabffabffab;
mem[5981] = 80'h0010ffabffabffabffab;
mem[5982] = 80'h0010ffabffabffabffab;
mem[5983] = 80'h0010ffabffabffabffab;
mem[5984] = 80'h0010ffabffabffabffab;
mem[5985] = 80'h0010ffabffabffabffab;
mem[5986] = 80'h0010ffabffabffabffab;
mem[5987] = 80'h0010ffabffabffabffab;
mem[5988] = 80'h0010ffabffabffabffab;
mem[5989] = 80'h0010ffabffabffabffab;
mem[5990] = 80'h0010ffabffabffabffab;
mem[5991] = 80'h0010ffabffabffabffab;
mem[5992] = 80'h0010ffabffabffabffab;
mem[5993] = 80'h0010ffabffabffabffab;
mem[5994] = 80'h0010ffabffabffabffab;
mem[5995] = 80'h0010ffabffabffabffab;
mem[5996] = 80'h0010ffabffabffabffab;
mem[5997] = 80'h0010ffabffabffabffab;
mem[5998] = 80'h0010ffabffabffabffab;
mem[5999] = 80'h0010ffabffabffabffab;
mem[6000] = 80'h0010ffabffabffabffab;
mem[6001] = 80'h0010ffabffabffabffab;
mem[6002] = 80'h0010ffabffabffabffab;
mem[6003] = 80'h0010ffabffabffabffab;
mem[6004] = 80'h0010ffabffabffabffab;
mem[6005] = 80'h0010ffabffabffabffab;
mem[6006] = 80'h0010ffabffabffabffab;
mem[6007] = 80'h0010ffabffabffabffab;
mem[6008] = 80'h0010ffabffabffabffab;
mem[6009] = 80'h0010ffabffabffabffab;
mem[6010] = 80'h0010ffabffabffabffab;
mem[6011] = 80'h0010ffabffabffabffab;
mem[6012] = 80'h0010ffabffabffabffab;
mem[6013] = 80'h0010ffabffabffabffab;
mem[6014] = 80'h0010ffabffabffabffab;
mem[6015] = 80'h0010ffabffabff2cd878;
mem[6016] = 80'h0010c2bf425af09a7c03;
mem[6017] = 80'h0010a0bdf934fed81bd7;
mem[6018] = 80'h011501a00edbf2000000;
mem[6019] = 80'h10100000010000010010;
mem[6020] = 80'h00109400000208004500;
mem[6021] = 80'h001003b189d40000fffd;
mem[6022] = 80'h0010ac22c0550102c000;
mem[6023] = 80'h00100001ffabffabffab;
mem[6024] = 80'h0010ffabffabffabffab;
mem[6025] = 80'h0010ffabffabffabffab;
mem[6026] = 80'h0010ffabffabffabffab;
mem[6027] = 80'h0010ffabffabffabffab;
mem[6028] = 80'h0010ffabffabffabffab;
mem[6029] = 80'h0010ffabffabffabffab;
mem[6030] = 80'h0010ffabffabffabffab;
mem[6031] = 80'h0010ffabffabffabffab;
mem[6032] = 80'h0010ffabffabffabffab;
mem[6033] = 80'h0010ffabffabffabffab;
mem[6034] = 80'h0010ffabffabffabffab;
mem[6035] = 80'h0010ffabffabffabffab;
mem[6036] = 80'h0010ffabffabffabffab;
mem[6037] = 80'h0010ffabffabffabffab;
mem[6038] = 80'h0010ffabffabffabffab;
mem[6039] = 80'h0010ffabffabffabffab;
mem[6040] = 80'h0010ffabffabffabffab;
mem[6041] = 80'h0010ffabffabffabffab;
mem[6042] = 80'h0010ffabffabffabffab;
mem[6043] = 80'h0010ffabffabffabffab;
mem[6044] = 80'h0010ffabffabffabffab;
mem[6045] = 80'h0010ffabffabffabffab;
mem[6046] = 80'h0010ffabffabffabffab;
mem[6047] = 80'h0010ffabffabffabffab;
mem[6048] = 80'h0010ffabffabffabffab;
mem[6049] = 80'h0010ffabffabffabffab;
mem[6050] = 80'h0010ffabffabffabffab;
mem[6051] = 80'h0010ffabffabffabffab;
mem[6052] = 80'h0010ffabffabffabffab;
mem[6053] = 80'h0010ffabffabffabffab;
mem[6054] = 80'h0010ffabffabffabffab;
mem[6055] = 80'h0010ffabffabffabffab;
mem[6056] = 80'h0010ffabffabffabffab;
mem[6057] = 80'h0010ffabffabffabffab;
mem[6058] = 80'h0010ffabffabffabffab;
mem[6059] = 80'h0010ffabffabffabffab;
mem[6060] = 80'h0010ffabffabffabffab;
mem[6061] = 80'h0010ffabffabffabffab;
mem[6062] = 80'h0010ffabffabffabffab;
mem[6063] = 80'h0010ffabffabffabffab;
mem[6064] = 80'h0010ffabffabffabffab;
mem[6065] = 80'h0010ffabffabffabffab;
mem[6066] = 80'h0010ffabffabffabffab;
mem[6067] = 80'h0010ffabffabffabffab;
mem[6068] = 80'h0010ffabffabffabffab;
mem[6069] = 80'h0010ffabffabffabffab;
mem[6070] = 80'h0010ffabffabffabffab;
mem[6071] = 80'h0010ffabffabffabffab;
mem[6072] = 80'h0010ffabffabffabffab;
mem[6073] = 80'h0010ffabffabffabffab;
mem[6074] = 80'h0010ffabffabffabffab;
mem[6075] = 80'h0010ffabffabffabffab;
mem[6076] = 80'h0010ffabffabffabffab;
mem[6077] = 80'h0010ffabffabffabffab;
mem[6078] = 80'h0010ffabffabffabffab;
mem[6079] = 80'h0010ffabffabffabffab;
mem[6080] = 80'h0010ffabffabffabffab;
mem[6081] = 80'h0010ffabffabffabffab;
mem[6082] = 80'h0010ffabffabffabffab;
mem[6083] = 80'h0010ffabffabffabffab;
mem[6084] = 80'h0010ffabffabffabffab;
mem[6085] = 80'h0010ffabffabffabffab;
mem[6086] = 80'h0010ffabffabffabffab;
mem[6087] = 80'h0010ffabffabffabffab;
mem[6088] = 80'h0010ffabffabffabffab;
mem[6089] = 80'h0010ffabffabffabffab;
mem[6090] = 80'h0010ffabffabffabffab;
mem[6091] = 80'h0010ffabffabffabffab;
mem[6092] = 80'h0010ffabffabffabffab;
mem[6093] = 80'h0010ffabffabffabffab;
mem[6094] = 80'h0010ffabffabffabffab;
mem[6095] = 80'h0010ffabffabffabffab;
mem[6096] = 80'h0010ffabffabffabffab;
mem[6097] = 80'h0010ffabffabffabffab;
mem[6098] = 80'h0010ffabffabffabffab;
mem[6099] = 80'h0010ffabffabffabffab;
mem[6100] = 80'h0010ffabffabffabffab;
mem[6101] = 80'h0010ffabffabffabffab;
mem[6102] = 80'h0010ffabffabffabffab;
mem[6103] = 80'h0010ffabffabffabffab;
mem[6104] = 80'h0010ffabffabffabffab;
mem[6105] = 80'h0010ffabffabffabffab;
mem[6106] = 80'h0010ffabffabffabffab;
mem[6107] = 80'h0010ffabffabffabffab;
mem[6108] = 80'h0010ffabffabffabffab;
mem[6109] = 80'h0010ffabffabffabffab;
mem[6110] = 80'h0010ffabffabffabffab;
mem[6111] = 80'h0010ffabffabffabffab;
mem[6112] = 80'h0010ffabffabffabffab;
mem[6113] = 80'h0010ffabffabffabffab;
mem[6114] = 80'h0010ffabffabffabffab;
mem[6115] = 80'h0010ffabffabffabffab;
mem[6116] = 80'h0010ffabffabffabffab;
mem[6117] = 80'h0010ffabffabffabffab;
mem[6118] = 80'h0010ffabffabffabffab;
mem[6119] = 80'h0010ffabffabffabffab;
mem[6120] = 80'h0010ffabffabffabffab;
mem[6121] = 80'h0010ffabffabffabffab;
mem[6122] = 80'h0010ffabffabffabffab;
mem[6123] = 80'h0010ffabffabffabffab;
mem[6124] = 80'h0010ffabffabffabffab;
mem[6125] = 80'h0010ffabffabffabffab;
mem[6126] = 80'h0010ffabffabffabffab;
mem[6127] = 80'h0010ffabffabffabffab;
mem[6128] = 80'h0010ffabffabffabffab;
mem[6129] = 80'h0010ffabffabffabffab;
mem[6130] = 80'h0010ffabffabffabffab;
mem[6131] = 80'h0010ffabffabffabffab;
mem[6132] = 80'h0010ffabffabffabffab;
mem[6133] = 80'h0010ffabffabffabffab;
mem[6134] = 80'h0010ffabffabffabffab;
mem[6135] = 80'h0010ffabffabffabffab;
mem[6136] = 80'h0010ffabff2bfcbc286e;
mem[6137] = 80'h001056d570229312cc81;
mem[6138] = 80'h001018e11b7796c4e99c;
mem[6139] = 80'h011395d3070000000000;
mem[6140] = 80'h10100000010000010010;
mem[6141] = 80'h00109400000208004500;
mem[6142] = 80'h001001ef89d50000fffd;
mem[6143] = 80'h0010ade3c0550102c000;
mem[6144] = 80'h00100001ffabffabffab;
mem[6145] = 80'h0010ffabffabffabffab;
mem[6146] = 80'h0010ffabffabffabffab;
mem[6147] = 80'h0010ffabffabffabffab;
mem[6148] = 80'h0010ffabffabffabffab;
mem[6149] = 80'h0010ffabffabffabffab;
mem[6150] = 80'h0010ffabffabffabffab;
mem[6151] = 80'h0010ffabffabffabffab;
mem[6152] = 80'h0010ffabffabffabffab;
mem[6153] = 80'h0010ffabffabffabffab;
mem[6154] = 80'h0010ffabffabffabffab;
mem[6155] = 80'h0010ffabffabffabffab;
mem[6156] = 80'h0010ffabffabffabffab;
mem[6157] = 80'h0010ffabffabffabffab;
mem[6158] = 80'h0010ffabffabffabffab;
mem[6159] = 80'h0010ffabffabffabffab;
mem[6160] = 80'h0010ffabffabffabffab;
mem[6161] = 80'h0010ffabffabffabffab;
mem[6162] = 80'h0010ffabffabffabffab;
mem[6163] = 80'h0010ffabffabffabffab;
mem[6164] = 80'h0010ffabffabffabffab;
mem[6165] = 80'h0010ffabffabffabffab;
mem[6166] = 80'h0010ffabffabffabffab;
mem[6167] = 80'h0010ffabffabffabffab;
mem[6168] = 80'h0010ffabffabffabffab;
mem[6169] = 80'h0010ffabffabffabffab;
mem[6170] = 80'h0010ffabffabffabffab;
mem[6171] = 80'h0010ffabffabffabffab;
mem[6172] = 80'h0010ffabffabffabffab;
mem[6173] = 80'h0010ffabffabffabffab;
mem[6174] = 80'h0010ffabffabffabffab;
mem[6175] = 80'h0010ffabffabffabffab;
mem[6176] = 80'h0010ffabffabffabffab;
mem[6177] = 80'h0010ffabffabffabffab;
mem[6178] = 80'h0010ffabffabffabffab;
mem[6179] = 80'h0010ffabffabffabffab;
mem[6180] = 80'h0010ffabffabffabffab;
mem[6181] = 80'h0010ffabffabffabffab;
mem[6182] = 80'h0010ffabffabffabffab;
mem[6183] = 80'h0010ffabffabffabffab;
mem[6184] = 80'h0010ffabffabffabffab;
mem[6185] = 80'h0010ffabffabffabffab;
mem[6186] = 80'h0010ffabffabffabffab;
mem[6187] = 80'h0010ffabffabffabffab;
mem[6188] = 80'h0010ffabffabffabffab;
mem[6189] = 80'h0010ffabffabffabffab;
mem[6190] = 80'h0010ffabffabffabffab;
mem[6191] = 80'h0010ffabffabffabffab;
mem[6192] = 80'h0010ffabffabffabffab;
mem[6193] = 80'h0010ffabffabffabffab;
mem[6194] = 80'h0010ffabffabffabffab;
mem[6195] = 80'h0010ffabffabffabffab;
mem[6196] = 80'h0010ffabffabffabffab;
mem[6197] = 80'h0010ffabffabffabffab;
mem[6198] = 80'h0010ffabffabffabffab;
mem[6199] = 80'h0010ffabffabffabffab;
mem[6200] = 80'h0010ffabffabffabffab;
mem[6201] = 80'h0010ff2a8d6204b62f17;
mem[6202] = 80'h0010cfe941952174ca43;
mem[6203] = 80'h00104a13205bd7054034;
mem[6204] = 80'h0111f100000000000000;
mem[6205] = 80'h10100000010000010010;
mem[6206] = 80'h00109400000208004500;
mem[6207] = 80'h0010011089d60000fffd;
mem[6208] = 80'h0010aec1c0550102c000;
mem[6209] = 80'h00100001ffabffabffab;
mem[6210] = 80'h0010ffabffabffabffab;
mem[6211] = 80'h0010ffabffabffabffab;
mem[6212] = 80'h0010ffabffabffabffab;
mem[6213] = 80'h0010ffabffabffabffab;
mem[6214] = 80'h0010ffabffabffabffab;
mem[6215] = 80'h0010ffabffabffabffab;
mem[6216] = 80'h0010ffabffabffabffab;
mem[6217] = 80'h0010ffabffabffabffab;
mem[6218] = 80'h0010ffabffabffabffab;
mem[6219] = 80'h0010ffabffabffabffab;
mem[6220] = 80'h0010ffabffabffabffab;
mem[6221] = 80'h0010ffabffabffabffab;
mem[6222] = 80'h0010ffabffabffabffab;
mem[6223] = 80'h0010ffabffabffabffab;
mem[6224] = 80'h0010ffabffabffabffab;
mem[6225] = 80'h0010ffabffabffabffab;
mem[6226] = 80'h0010ffabffabffabffab;
mem[6227] = 80'h0010ffabffabffabffab;
mem[6228] = 80'h0010ffabffabffabffab;
mem[6229] = 80'h0010ffabffabffabffab;
mem[6230] = 80'h0010ffabffabffabffab;
mem[6231] = 80'h0010ffabffabffabffab;
mem[6232] = 80'h0010ffabffabffabffab;
mem[6233] = 80'h0010ffabffabffabffab;
mem[6234] = 80'h0010ffabffabffabffab;
mem[6235] = 80'h0010ffabffabffabffab;
mem[6236] = 80'h0010ffabffabffabffab;
mem[6237] = 80'h0010ffabffabffabffab;
mem[6238] = 80'h0010ffab291f0071dea5;
mem[6239] = 80'h0010500fb5361d176aba;
mem[6240] = 80'h001031b8ff643995be15;
mem[6241] = 80'h0112a9fa000000000000;
mem[6242] = 80'h10100000010000010010;
mem[6243] = 80'h00109400000208004500;
mem[6244] = 80'h0010009f89d70000fffd;
mem[6245] = 80'h0010af31c0550102c000;
mem[6246] = 80'h00100001ffabffabffab;
mem[6247] = 80'h0010ffabffabffabffab;
mem[6248] = 80'h0010ffabffabffabffab;
mem[6249] = 80'h0010ffabffabffabffab;
mem[6250] = 80'h0010ffabffabffabffab;
mem[6251] = 80'h0010ffabffabffabffab;
mem[6252] = 80'h0010ffabffabffabffab;
mem[6253] = 80'h0010ffabffabffabffab;
mem[6254] = 80'h0010ffabffabffabffab;
mem[6255] = 80'h0010ffabffabffabffab;
mem[6256] = 80'h0010ffabffabffabffab;
mem[6257] = 80'h0010ffabffabffabffab;
mem[6258] = 80'h0010ffabffabffabffab;
mem[6259] = 80'h0010ffabffabffabffab;
mem[6260] = 80'h0010ffabffabffabffab;
mem[6261] = 80'h0010ff286ede5d06dc92;
mem[6262] = 80'h0010b07ee49afa9f65b8;
mem[6263] = 80'h0010e9039fe9d9d2f863;
mem[6264] = 80'h01113800000000000000;
mem[6265] = 80'h10100000010000010010;
mem[6266] = 80'h00109400000208004500;
mem[6267] = 80'h0010006589d80000fffd;
mem[6268] = 80'h0010af6ac0550102c000;
mem[6269] = 80'h00100001ffabffabffab;
mem[6270] = 80'h0010ffabffabffabffab;
mem[6271] = 80'h0010ffabffabffabffab;
mem[6272] = 80'h0010ffabffabffabffab;
mem[6273] = 80'h0010ffabffabffabffab;
mem[6274] = 80'h0010ffabffabffabffab;
mem[6275] = 80'h0010ffabffabffabffab;
mem[6276] = 80'h0010ffabffabffabff27;
mem[6277] = 80'h00105689a47c8c4f0ec4;
mem[6278] = 80'h0010e83fcf137722732c;
mem[6279] = 80'h0117db1bed1dc721e600;
mem[6280] = 80'h10100000010000010010;
mem[6281] = 80'h00109400000208004500;
mem[6282] = 80'h0010032189d90000fffd;
mem[6283] = 80'h0010acadc0550102c000;
mem[6284] = 80'h00100001ffabffabffab;
mem[6285] = 80'h0010ffabffabffabffab;
mem[6286] = 80'h0010ffabffabffabffab;
mem[6287] = 80'h0010ffabffabffabffab;
mem[6288] = 80'h0010ffabffabffabffab;
mem[6289] = 80'h0010ffabffabffabffab;
mem[6290] = 80'h0010ffabffabffabffab;
mem[6291] = 80'h0010ffabffabffabffab;
mem[6292] = 80'h0010ffabffabffabffab;
mem[6293] = 80'h0010ffabffabffabffab;
mem[6294] = 80'h0010ffabffabffabffab;
mem[6295] = 80'h0010ffabffabffabffab;
mem[6296] = 80'h0010ffabffabffabffab;
mem[6297] = 80'h0010ffabffabffabffab;
mem[6298] = 80'h0010ffabffabffabffab;
mem[6299] = 80'h0010ffabffabffabffab;
mem[6300] = 80'h0010ffabffabffabffab;
mem[6301] = 80'h0010ffabffabffabffab;
mem[6302] = 80'h0010ffabffabffabffab;
mem[6303] = 80'h0010ffabffabffabffab;
mem[6304] = 80'h0010ffabffabffabffab;
mem[6305] = 80'h0010ffabffabffabffab;
mem[6306] = 80'h0010ffabffabffabffab;
mem[6307] = 80'h0010ffabffabffabffab;
mem[6308] = 80'h0010ffabffabffabffab;
mem[6309] = 80'h0010ffabffabffabffab;
mem[6310] = 80'h0010ffabffabffabffab;
mem[6311] = 80'h0010ffabffabffabffab;
mem[6312] = 80'h0010ffabffabffabffab;
mem[6313] = 80'h0010ffabffabffabffab;
mem[6314] = 80'h0010ffabffabffabffab;
mem[6315] = 80'h0010ffabffabffabffab;
mem[6316] = 80'h0010ffabffabffabffab;
mem[6317] = 80'h0010ffabffabffabffab;
mem[6318] = 80'h0010ffabffabffabffab;
mem[6319] = 80'h0010ffabffabffabffab;
mem[6320] = 80'h0010ffabffabffabffab;
mem[6321] = 80'h0010ffabffabffabffab;
mem[6322] = 80'h0010ffabffabffabffab;
mem[6323] = 80'h0010ffabffabffabffab;
mem[6324] = 80'h0010ffabffabffabffab;
mem[6325] = 80'h0010ffabffabffabffab;
mem[6326] = 80'h0010ffabffabffabffab;
mem[6327] = 80'h0010ffabffabffabffab;
mem[6328] = 80'h0010ffabffabffabffab;
mem[6329] = 80'h0010ffabffabffabffab;
mem[6330] = 80'h0010ffabffabffabffab;
mem[6331] = 80'h0010ffabffabffabffab;
mem[6332] = 80'h0010ffabffabffabffab;
mem[6333] = 80'h0010ffabffabffabffab;
mem[6334] = 80'h0010ffabffabffabffab;
mem[6335] = 80'h0010ffabffabffabffab;
mem[6336] = 80'h0010ffabffabffabffab;
mem[6337] = 80'h0010ffabffabffabffab;
mem[6338] = 80'h0010ffabffabffabffab;
mem[6339] = 80'h0010ffabffabffabffab;
mem[6340] = 80'h0010ffabffabffabffab;
mem[6341] = 80'h0010ffabffabffabffab;
mem[6342] = 80'h0010ffabffabffabffab;
mem[6343] = 80'h0010ffabffabffabffab;
mem[6344] = 80'h0010ffabffabffabffab;
mem[6345] = 80'h0010ffabffabffabffab;
mem[6346] = 80'h0010ffabffabffabffab;
mem[6347] = 80'h0010ffabffabffabffab;
mem[6348] = 80'h0010ffabffabffabffab;
mem[6349] = 80'h0010ffabffabffabffab;
mem[6350] = 80'h0010ffabffabffabffab;
mem[6351] = 80'h0010ffabffabffabffab;
mem[6352] = 80'h0010ffabffabffabffab;
mem[6353] = 80'h0010ffabffabffabffab;
mem[6354] = 80'h0010ffabffabffabffab;
mem[6355] = 80'h0010ffabffabffabffab;
mem[6356] = 80'h0010ffabffabffabffab;
mem[6357] = 80'h0010ffabffabffabffab;
mem[6358] = 80'h0010ffabffabffabffab;
mem[6359] = 80'h0010ffabffabffabffab;
mem[6360] = 80'h0010ffabffabffabffab;
mem[6361] = 80'h0010ffabffabffabffab;
mem[6362] = 80'h0010ffabffabffabffab;
mem[6363] = 80'h0010ffabffabffabffab;
mem[6364] = 80'h0010ffabffabffabffab;
mem[6365] = 80'h0010ffabffabffabffab;
mem[6366] = 80'h0010ffabffabffabffab;
mem[6367] = 80'h0010ffabffabffabffab;
mem[6368] = 80'h0010ffabffabffabffab;
mem[6369] = 80'h0010ffabffabffabffab;
mem[6370] = 80'h0010ffabffabffabffab;
mem[6371] = 80'h0010ffabffabffabffab;
mem[6372] = 80'h0010ffabffabffabffab;
mem[6373] = 80'h0010ffabffabffabffab;
mem[6374] = 80'h0010ffabffabffabffab;
mem[6375] = 80'h0010ffabffabffabffab;
mem[6376] = 80'h0010ffabffabffabffab;
mem[6377] = 80'h0010ffabffabffabffab;
mem[6378] = 80'h0010ffabffabffabffab;
mem[6379] = 80'h0010ffabff26275788a4;
mem[6380] = 80'h0010f58db10f3ab822e6;
mem[6381] = 80'h0010a7bb22ff62e71e9b;
mem[6382] = 80'h0113683dee0000000000;
mem[6383] = 80'h10100000010000010010;
mem[6384] = 80'h00109400000208004500;
mem[6385] = 80'h0010047d89da0000fffd;
mem[6386] = 80'h0010ab50c0550102c000;
mem[6387] = 80'h00100001ffabffabffab;
mem[6388] = 80'h0010ffabffabffabffab;
mem[6389] = 80'h0010ffabffabffabffab;
mem[6390] = 80'h0010ffabffabffabffab;
mem[6391] = 80'h0010ffabffabffabffab;
mem[6392] = 80'h0010ffabffabffabffab;
mem[6393] = 80'h0010ffabffabffabffab;
mem[6394] = 80'h0010ffabffabffabffab;
mem[6395] = 80'h0010ffabffabffabffab;
mem[6396] = 80'h0010ffabffabffabffab;
mem[6397] = 80'h0010ffabffabffabffab;
mem[6398] = 80'h0010ffabffabffabffab;
mem[6399] = 80'h0010ffabffabffabffab;
mem[6400] = 80'h0010ffabffabffabffab;
mem[6401] = 80'h0010ffabffabffabffab;
mem[6402] = 80'h0010ffabffabffabffab;
mem[6403] = 80'h0010ffabffabffabffab;
mem[6404] = 80'h0010ffabffabffabffab;
mem[6405] = 80'h0010ffabffabffabffab;
mem[6406] = 80'h0010ffabffabffabffab;
mem[6407] = 80'h0010ffabffabffabffab;
mem[6408] = 80'h0010ffabffabffabffab;
mem[6409] = 80'h0010ffabffabffabffab;
mem[6410] = 80'h0010ffabffabffabffab;
mem[6411] = 80'h0010ffabffabffabffab;
mem[6412] = 80'h0010ffabffabffabffab;
mem[6413] = 80'h0010ffabffabffabffab;
mem[6414] = 80'h0010ffabffabffabffab;
mem[6415] = 80'h0010ffabffabffabffab;
mem[6416] = 80'h0010ffabffabffabffab;
mem[6417] = 80'h0010ffabffabffabffab;
mem[6418] = 80'h0010ffabffabffabffab;
mem[6419] = 80'h0010ffabffabffabffab;
mem[6420] = 80'h0010ffabffabffabffab;
mem[6421] = 80'h0010ffabffabffabffab;
mem[6422] = 80'h0010ffabffabffabffab;
mem[6423] = 80'h0010ffabffabffabffab;
mem[6424] = 80'h0010ffabffabffabffab;
mem[6425] = 80'h0010ffabffabffabffab;
mem[6426] = 80'h0010ffabffabffabffab;
mem[6427] = 80'h0010ffabffabffabffab;
mem[6428] = 80'h0010ffabffabffabffab;
mem[6429] = 80'h0010ffabffabffabffab;
mem[6430] = 80'h0010ffabffabffabffab;
mem[6431] = 80'h0010ffabffabffabffab;
mem[6432] = 80'h0010ffabffabffabffab;
mem[6433] = 80'h0010ffabffabffabffab;
mem[6434] = 80'h0010ffabffabffabffab;
mem[6435] = 80'h0010ffabffabffabffab;
mem[6436] = 80'h0010ffabffabffabffab;
mem[6437] = 80'h0010ffabffabffabffab;
mem[6438] = 80'h0010ffabffabffabffab;
mem[6439] = 80'h0010ffabffabffabffab;
mem[6440] = 80'h0010ffabffabffabffab;
mem[6441] = 80'h0010ffabffabffabffab;
mem[6442] = 80'h0010ffabffabffabffab;
mem[6443] = 80'h0010ffabffabffabffab;
mem[6444] = 80'h0010ffabffabffabffab;
mem[6445] = 80'h0010ffabffabffabffab;
mem[6446] = 80'h0010ffabffabffabffab;
mem[6447] = 80'h0010ffabffabffabffab;
mem[6448] = 80'h0010ffabffabffabffab;
mem[6449] = 80'h0010ffabffabffabffab;
mem[6450] = 80'h0010ffabffabffabffab;
mem[6451] = 80'h0010ffabffabffabffab;
mem[6452] = 80'h0010ffabffabffabffab;
mem[6453] = 80'h0010ffabffabffabffab;
mem[6454] = 80'h0010ffabffabffabffab;
mem[6455] = 80'h0010ffabffabffabffab;
mem[6456] = 80'h0010ffabffabffabffab;
mem[6457] = 80'h0010ffabffabffabffab;
mem[6458] = 80'h0010ffabffabffabffab;
mem[6459] = 80'h0010ffabffabffabffab;
mem[6460] = 80'h0010ffabffabffabffab;
mem[6461] = 80'h0010ffabffabffabffab;
mem[6462] = 80'h0010ffabffabffabffab;
mem[6463] = 80'h0010ffabffabffabffab;
mem[6464] = 80'h0010ffabffabffabffab;
mem[6465] = 80'h0010ffabffabffabffab;
mem[6466] = 80'h0010ffabffabffabffab;
mem[6467] = 80'h0010ffabffabffabffab;
mem[6468] = 80'h0010ffabffabffabffab;
mem[6469] = 80'h0010ffabffabffabffab;
mem[6470] = 80'h0010ffabffabffabffab;
mem[6471] = 80'h0010ffabffabffabffab;
mem[6472] = 80'h0010ffabffabffabffab;
mem[6473] = 80'h0010ffabffabffabffab;
mem[6474] = 80'h0010ffabffabffabffab;
mem[6475] = 80'h0010ffabffabffabffab;
mem[6476] = 80'h0010ffabffabffabffab;
mem[6477] = 80'h0010ffabffabffabffab;
mem[6478] = 80'h0010ffabffabffabffab;
mem[6479] = 80'h0010ffabffabffabffab;
mem[6480] = 80'h0010ffabffabffabffab;
mem[6481] = 80'h0010ffabffabffabffab;
mem[6482] = 80'h0010ffabffabffabffab;
mem[6483] = 80'h0010ffabffabffabffab;
mem[6484] = 80'h0010ffabffabffabffab;
mem[6485] = 80'h0010ffabffabffabffab;
mem[6486] = 80'h0010ffabffabffabffab;
mem[6487] = 80'h0010ffabffabffabffab;
mem[6488] = 80'h0010ffabffabffabffab;
mem[6489] = 80'h0010ffabffabffabffab;
mem[6490] = 80'h0010ffabffabffabffab;
mem[6491] = 80'h0010ffabffabffabffab;
mem[6492] = 80'h0010ffabffabffabffab;
mem[6493] = 80'h0010ffabffabffabffab;
mem[6494] = 80'h0010ffabffabffabffab;
mem[6495] = 80'h0010ffabffabffabffab;
mem[6496] = 80'h0010ffabffabffabffab;
mem[6497] = 80'h0010ffabffabffabffab;
mem[6498] = 80'h0010ffabffabffabffab;
mem[6499] = 80'h0010ffabffabffabffab;
mem[6500] = 80'h0010ffabffabffabffab;
mem[6501] = 80'h0010ffabffabffabffab;
mem[6502] = 80'h0010ffabffabffabffab;
mem[6503] = 80'h0010ffabffabffabffab;
mem[6504] = 80'h0010ffabffabffabffab;
mem[6505] = 80'h0010ffabffabffabffab;
mem[6506] = 80'h0010ffabffabffabffab;
mem[6507] = 80'h0010ffabffabffabffab;
mem[6508] = 80'h0010ffabffabffabffab;
mem[6509] = 80'h0010ffabffabffabffab;
mem[6510] = 80'h0010ffabffabffabffab;
mem[6511] = 80'h0010ffabffabffabffab;
mem[6512] = 80'h0010ffabffabffabffab;
mem[6513] = 80'h0010ffabffabffabffab;
mem[6514] = 80'h0010ffabffabffabffab;
mem[6515] = 80'h0010ffabffabffabffab;
mem[6516] = 80'h0010ffabffabffabffab;
mem[6517] = 80'h0010ffabffabffabffab;
mem[6518] = 80'h0010ffabffabffabffab;
mem[6519] = 80'h0010ffabffabffabffab;
mem[6520] = 80'h0010ffabffabffabffab;
mem[6521] = 80'h0010ffabffabffabffab;
mem[6522] = 80'h0010ffabffabffabffab;
mem[6523] = 80'h0010ffabffabffabffab;
mem[6524] = 80'h0010ffabffabffabffab;
mem[6525] = 80'h0010ffabffabffabff25;
mem[6526] = 80'h0010b535fdcc7fca7153;
mem[6527] = 80'h00104d3014f8d621d0bd;
mem[6528] = 80'h01170db2455466d46800;
mem[6529] = 80'h10100000010000010010;
mem[6530] = 80'h00109400000208004500;
mem[6531] = 80'h0010025589db0000fffd;
mem[6532] = 80'h0010ad77c0550102c000;
mem[6533] = 80'h00100001ffabffabffab;
mem[6534] = 80'h0010ffabffabffabffab;
mem[6535] = 80'h0010ffabffabffabffab;
mem[6536] = 80'h0010ffabffabffabffab;
mem[6537] = 80'h0010ffabffabffabffab;
mem[6538] = 80'h0010ffabffabffabffab;
mem[6539] = 80'h0010ffabffabffabffab;
mem[6540] = 80'h0010ffabffabffabffab;
mem[6541] = 80'h0010ffabffabffabffab;
mem[6542] = 80'h0010ffabffabffabffab;
mem[6543] = 80'h0010ffabffabffabffab;
mem[6544] = 80'h0010ffabffabffabffab;
mem[6545] = 80'h0010ffabffabffabffab;
mem[6546] = 80'h0010ffabffabffabffab;
mem[6547] = 80'h0010ffabffabffabffab;
mem[6548] = 80'h0010ffabffabffabffab;
mem[6549] = 80'h0010ffabffabffabffab;
mem[6550] = 80'h0010ffabffabffabffab;
mem[6551] = 80'h0010ffabffabffabffab;
mem[6552] = 80'h0010ffabffabffabffab;
mem[6553] = 80'h0010ffabffabffabffab;
mem[6554] = 80'h0010ffabffabffabffab;
mem[6555] = 80'h0010ffabffabffabffab;
mem[6556] = 80'h0010ffabffabffabffab;
mem[6557] = 80'h0010ffabffabffabffab;
mem[6558] = 80'h0010ffabffabffabffab;
mem[6559] = 80'h0010ffabffabffabffab;
mem[6560] = 80'h0010ffabffabffabffab;
mem[6561] = 80'h0010ffabffabffabffab;
mem[6562] = 80'h0010ffabffabffabffab;
mem[6563] = 80'h0010ffabffabffabffab;
mem[6564] = 80'h0010ffabffabffabffab;
mem[6565] = 80'h0010ffabffabffabffab;
mem[6566] = 80'h0010ffabffabffabffab;
mem[6567] = 80'h0010ffabffabffabffab;
mem[6568] = 80'h0010ffabffabffabffab;
mem[6569] = 80'h0010ffabffabffabffab;
mem[6570] = 80'h0010ffabffabffabffab;
mem[6571] = 80'h0010ffabffabffabffab;
mem[6572] = 80'h0010ffabffabffabffab;
mem[6573] = 80'h0010ffabffabffabffab;
mem[6574] = 80'h0010ffabffabffabffab;
mem[6575] = 80'h0010ffabffabffabffab;
mem[6576] = 80'h0010ffabffabffabffab;
mem[6577] = 80'h0010ffabffabffabffab;
mem[6578] = 80'h0010ffabffabffabffab;
mem[6579] = 80'h0010ffabffabffabffab;
mem[6580] = 80'h0010ffabffabffabffab;
mem[6581] = 80'h0010ffabffabffabffab;
mem[6582] = 80'h0010ffabffabffabffab;
mem[6583] = 80'h0010ffabffabffabffab;
mem[6584] = 80'h0010ffabffabffabffab;
mem[6585] = 80'h0010ffabffabffabffab;
mem[6586] = 80'h0010ffabffabffabffab;
mem[6587] = 80'h0010ffabffabffabffab;
mem[6588] = 80'h0010ffabffabffabffab;
mem[6589] = 80'h0010ffabffabffabffab;
mem[6590] = 80'h0010ffabffabffabffab;
mem[6591] = 80'h0010ffabffabffabffab;
mem[6592] = 80'h0010ffabffabffabffab;
mem[6593] = 80'h0010ffabffabffabffab;
mem[6594] = 80'h0010ffabffabffabffab;
mem[6595] = 80'h0010ffabffabffabffab;
mem[6596] = 80'h0010ffabffabffabffab;
mem[6597] = 80'h0010ffabffabffabffab;
mem[6598] = 80'h0010ffabffabffabffab;
mem[6599] = 80'h0010ffabffabffabffab;
mem[6600] = 80'h0010ffabffabffabffab;
mem[6601] = 80'h0010ffabffabffabffab;
mem[6602] = 80'h0010ffabffabffabff24;
mem[6603] = 80'h0010c4ebd1140608ce98;
mem[6604] = 80'h00109fb7f90d04fb8158;
mem[6605] = 80'h01174b212b833a6c9c00;
mem[6606] = 80'h10100000010000010010;
mem[6607] = 80'h00109400000208004500;
mem[6608] = 80'h0010041a89dc0000fffd;
mem[6609] = 80'h0010abb1c0550102c000;
mem[6610] = 80'h00100001ffabffabffab;
mem[6611] = 80'h0010ffabffabffabffab;
mem[6612] = 80'h0010ffabffabffabffab;
mem[6613] = 80'h0010ffabffabffabffab;
mem[6614] = 80'h0010ffabffabffabffab;
mem[6615] = 80'h0010ffabffabffabffab;
mem[6616] = 80'h0010ffabffabffabffab;
mem[6617] = 80'h0010ffabffabffabffab;
mem[6618] = 80'h0010ffabffabffabffab;
mem[6619] = 80'h0010ffabffabffabffab;
mem[6620] = 80'h0010ffabffabffabffab;
mem[6621] = 80'h0010ffabffabffabffab;
mem[6622] = 80'h0010ffabffabffabffab;
mem[6623] = 80'h0010ffabffabffabffab;
mem[6624] = 80'h0010ffabffabffabffab;
mem[6625] = 80'h0010ffabffabffabffab;
mem[6626] = 80'h0010ffabffabffabffab;
mem[6627] = 80'h0010ffabffabffabffab;
mem[6628] = 80'h0010ffabffabffabffab;
mem[6629] = 80'h0010ffabffabffabffab;
mem[6630] = 80'h0010ffabffabffabffab;
mem[6631] = 80'h0010ffabffabffabffab;
mem[6632] = 80'h0010ffabffabffabffab;
mem[6633] = 80'h0010ffabffabffabffab;
mem[6634] = 80'h0010ffabffabffabffab;
mem[6635] = 80'h0010ffabffabffabffab;
mem[6636] = 80'h0010ffabffabffabffab;
mem[6637] = 80'h0010ffabffabffabffab;
mem[6638] = 80'h0010ffabffabffabffab;
mem[6639] = 80'h0010ffabffabffabffab;
mem[6640] = 80'h0010ffabffabffabffab;
mem[6641] = 80'h0010ffabffabffabffab;
mem[6642] = 80'h0010ffabffabffabffab;
mem[6643] = 80'h0010ffabffabffabffab;
mem[6644] = 80'h0010ffabffabffabffab;
mem[6645] = 80'h0010ffabffabffabffab;
mem[6646] = 80'h0010ffabffabffabffab;
mem[6647] = 80'h0010ffabffabffabffab;
mem[6648] = 80'h0010ffabffabffabffab;
mem[6649] = 80'h0010ffabffabffabffab;
mem[6650] = 80'h0010ffabffabffabffab;
mem[6651] = 80'h0010ffabffabffabffab;
mem[6652] = 80'h0010ffabffabffabffab;
mem[6653] = 80'h0010ffabffabffabffab;
mem[6654] = 80'h0010ffabffabffabffab;
mem[6655] = 80'h0010ffabffabffabffab;
mem[6656] = 80'h0010ffabffabffabffab;
mem[6657] = 80'h0010ffabffabffabffab;
mem[6658] = 80'h0010ffabffabffabffab;
mem[6659] = 80'h0010ffabffabffabffab;
mem[6660] = 80'h0010ffabffabffabffab;
mem[6661] = 80'h0010ffabffabffabffab;
mem[6662] = 80'h0010ffabffabffabffab;
mem[6663] = 80'h0010ffabffabffabffab;
mem[6664] = 80'h0010ffabffabffabffab;
mem[6665] = 80'h0010ffabffabffabffab;
mem[6666] = 80'h0010ffabffabffabffab;
mem[6667] = 80'h0010ffabffabffabffab;
mem[6668] = 80'h0010ffabffabffabffab;
mem[6669] = 80'h0010ffabffabffabffab;
mem[6670] = 80'h0010ffabffabffabffab;
mem[6671] = 80'h0010ffabffabffabffab;
mem[6672] = 80'h0010ffabffabffabffab;
mem[6673] = 80'h0010ffabffabffabffab;
mem[6674] = 80'h0010ffabffabffabffab;
mem[6675] = 80'h0010ffabffabffabffab;
mem[6676] = 80'h0010ffabffabffabffab;
mem[6677] = 80'h0010ffabffabffabffab;
mem[6678] = 80'h0010ffabffabffabffab;
mem[6679] = 80'h0010ffabffabffabffab;
mem[6680] = 80'h0010ffabffabffabffab;
mem[6681] = 80'h0010ffabffabffabffab;
mem[6682] = 80'h0010ffabffabffabffab;
mem[6683] = 80'h0010ffabffabffabffab;
mem[6684] = 80'h0010ffabffabffabffab;
mem[6685] = 80'h0010ffabffabffabffab;
mem[6686] = 80'h0010ffabffabffabffab;
mem[6687] = 80'h0010ffabffabffabffab;
mem[6688] = 80'h0010ffabffabffabffab;
mem[6689] = 80'h0010ffabffabffabffab;
mem[6690] = 80'h0010ffabffabffabffab;
mem[6691] = 80'h0010ffabffabffabffab;
mem[6692] = 80'h0010ffabffabffabffab;
mem[6693] = 80'h0010ffabffabffabffab;
mem[6694] = 80'h0010ffabffabffabffab;
mem[6695] = 80'h0010ffabffabffabffab;
mem[6696] = 80'h0010ffabffabffabffab;
mem[6697] = 80'h0010ffabffabffabffab;
mem[6698] = 80'h0010ffabffabffabffab;
mem[6699] = 80'h0010ffabffabffabffab;
mem[6700] = 80'h0010ffabffabffabffab;
mem[6701] = 80'h0010ffabffabffabffab;
mem[6702] = 80'h0010ffabffabffabffab;
mem[6703] = 80'h0010ffabffabffabffab;
mem[6704] = 80'h0010ffabffabffabffab;
mem[6705] = 80'h0010ffabffabffabffab;
mem[6706] = 80'h0010ffabffabffabffab;
mem[6707] = 80'h0010ffabffabffabffab;
mem[6708] = 80'h0010ffabffabffabffab;
mem[6709] = 80'h0010ffabffabffabffab;
mem[6710] = 80'h0010ffabffabffabffab;
mem[6711] = 80'h0010ffabffabffabffab;
mem[6712] = 80'h0010ffabffabffabffab;
mem[6713] = 80'h0010ffabffabffabffab;
mem[6714] = 80'h0010ffabffabffabffab;
mem[6715] = 80'h0010ffabffabffabffab;
mem[6716] = 80'h0010ffabffabffabffab;
mem[6717] = 80'h0010ffabffabffabffab;
mem[6718] = 80'h0010ffabffabffabffab;
mem[6719] = 80'h0010ffabffabffabffab;
mem[6720] = 80'h0010ffabffabffabffab;
mem[6721] = 80'h0010ffabffabffabffab;
mem[6722] = 80'h0010ffabffabffabffab;
mem[6723] = 80'h0010ffabffabffabffab;
mem[6724] = 80'h0010ffabffabffabffab;
mem[6725] = 80'h0010ffabffabffabffab;
mem[6726] = 80'h0010ffabffabffabffab;
mem[6727] = 80'h0010ffabffabffabffab;
mem[6728] = 80'h0010ffabffabffabffab;
mem[6729] = 80'h0010ffabffabffabffab;
mem[6730] = 80'h0010ffabffabffabffab;
mem[6731] = 80'h0010ffabffabffabffab;
mem[6732] = 80'h0010ffabffabffabffab;
mem[6733] = 80'h0010ffabffabffabffab;
mem[6734] = 80'h0010ffabffabffabffab;
mem[6735] = 80'h0010ffabffabffabffab;
mem[6736] = 80'h0010ffabffab23e02f3b;
mem[6737] = 80'h0010c512874e2070a695;
mem[6738] = 80'h001031e5536489c38a70;
mem[6739] = 80'h01146f5571a000000000;
mem[6740] = 80'h10100000010000010010;
mem[6741] = 80'h00109400000208004500;
mem[6742] = 80'h0010022489dd0000fffd;
mem[6743] = 80'h0010ada6c0550102c000;
mem[6744] = 80'h00100001ffabffabffab;
mem[6745] = 80'h0010ffabffabffabffab;
mem[6746] = 80'h0010ffabffabffabffab;
mem[6747] = 80'h0010ffabffabffabffab;
mem[6748] = 80'h0010ffabffabffabffab;
mem[6749] = 80'h0010ffabffabffabffab;
mem[6750] = 80'h0010ffabffabffabffab;
mem[6751] = 80'h0010ffabffabffabffab;
mem[6752] = 80'h0010ffabffabffabffab;
mem[6753] = 80'h0010ffabffabffabffab;
mem[6754] = 80'h0010ffabffabffabffab;
mem[6755] = 80'h0010ffabffabffabffab;
mem[6756] = 80'h0010ffabffabffabffab;
mem[6757] = 80'h0010ffabffabffabffab;
mem[6758] = 80'h0010ffabffabffabffab;
mem[6759] = 80'h0010ffabffabffabffab;
mem[6760] = 80'h0010ffabffabffabffab;
mem[6761] = 80'h0010ffabffabffabffab;
mem[6762] = 80'h0010ffabffabffabffab;
mem[6763] = 80'h0010ffabffabffabffab;
mem[6764] = 80'h0010ffabffabffabffab;
mem[6765] = 80'h0010ffabffabffabffab;
mem[6766] = 80'h0010ffabffabffabffab;
mem[6767] = 80'h0010ffabffabffabffab;
mem[6768] = 80'h0010ffabffabffabffab;
mem[6769] = 80'h0010ffabffabffabffab;
mem[6770] = 80'h0010ffabffabffabffab;
mem[6771] = 80'h0010ffabffabffabffab;
mem[6772] = 80'h0010ffabffabffabffab;
mem[6773] = 80'h0010ffabffabffabffab;
mem[6774] = 80'h0010ffabffabffabffab;
mem[6775] = 80'h0010ffabffabffabffab;
mem[6776] = 80'h0010ffabffabffabffab;
mem[6777] = 80'h0010ffabffabffabffab;
mem[6778] = 80'h0010ffabffabffabffab;
mem[6779] = 80'h0010ffabffabffabffab;
mem[6780] = 80'h0010ffabffabffabffab;
mem[6781] = 80'h0010ffabffabffabffab;
mem[6782] = 80'h0010ffabffabffabffab;
mem[6783] = 80'h0010ffabffabffabffab;
mem[6784] = 80'h0010ffabffabffabffab;
mem[6785] = 80'h0010ffabffabffabffab;
mem[6786] = 80'h0010ffabffabffabffab;
mem[6787] = 80'h0010ffabffabffabffab;
mem[6788] = 80'h0010ffabffabffabffab;
mem[6789] = 80'h0010ffabffabffabffab;
mem[6790] = 80'h0010ffabffabffabffab;
mem[6791] = 80'h0010ffabffabffabffab;
mem[6792] = 80'h0010ffabffabffabffab;
mem[6793] = 80'h0010ffabffabffabffab;
mem[6794] = 80'h0010ffabffabffabffab;
mem[6795] = 80'h0010ffabffabffabffab;
mem[6796] = 80'h0010ffabffabffabffab;
mem[6797] = 80'h0010ffabffabffabffab;
mem[6798] = 80'h0010ffabffabffabffab;
mem[6799] = 80'h0010ffabffabffabffab;
mem[6800] = 80'h0010ffabffabffabffab;
mem[6801] = 80'h0010ffabffabffabffab;
mem[6802] = 80'h0010ffabffabffabffab;
mem[6803] = 80'h0010ffabffabffabffab;
mem[6804] = 80'h0010ffabffabffabffab;
mem[6805] = 80'h0010ffabffabffabffab;
mem[6806] = 80'h0010ffabffabffabffab;
mem[6807] = 80'h0010ffabffabffab2291;
mem[6808] = 80'h0010f1171d6b45f1eba2;
mem[6809] = 80'h00102178c43398358007;
mem[6810] = 80'h01169f6ec266703d0000;
mem[6811] = 80'h10100000010000010010;
mem[6812] = 80'h00109400000208004500;
mem[6813] = 80'h0010040089de0000fffd;
mem[6814] = 80'h0010abc9c0550102c000;
mem[6815] = 80'h00100001ffabffabffab;
mem[6816] = 80'h0010ffabffabffabffab;
mem[6817] = 80'h0010ffabffabffabffab;
mem[6818] = 80'h0010ffabffabffabffab;
mem[6819] = 80'h0010ffabffabffabffab;
mem[6820] = 80'h0010ffabffabffabffab;
mem[6821] = 80'h0010ffabffabffabffab;
mem[6822] = 80'h0010ffabffabffabffab;
mem[6823] = 80'h0010ffabffabffabffab;
mem[6824] = 80'h0010ffabffabffabffab;
mem[6825] = 80'h0010ffabffabffabffab;
mem[6826] = 80'h0010ffabffabffabffab;
mem[6827] = 80'h0010ffabffabffabffab;
mem[6828] = 80'h0010ffabffabffabffab;
mem[6829] = 80'h0010ffabffabffabffab;
mem[6830] = 80'h0010ffabffabffabffab;
mem[6831] = 80'h0010ffabffabffabffab;
mem[6832] = 80'h0010ffabffabffabffab;
mem[6833] = 80'h0010ffabffabffabffab;
mem[6834] = 80'h0010ffabffabffabffab;
mem[6835] = 80'h0010ffabffabffabffab;
mem[6836] = 80'h0010ffabffabffabffab;
mem[6837] = 80'h0010ffabffabffabffab;
mem[6838] = 80'h0010ffabffabffabffab;
mem[6839] = 80'h0010ffabffabffabffab;
mem[6840] = 80'h0010ffabffabffabffab;
mem[6841] = 80'h0010ffabffabffabffab;
mem[6842] = 80'h0010ffabffabffabffab;
mem[6843] = 80'h0010ffabffabffabffab;
mem[6844] = 80'h0010ffabffabffabffab;
mem[6845] = 80'h0010ffabffabffabffab;
mem[6846] = 80'h0010ffabffabffabffab;
mem[6847] = 80'h0010ffabffabffabffab;
mem[6848] = 80'h0010ffabffabffabffab;
mem[6849] = 80'h0010ffabffabffabffab;
mem[6850] = 80'h0010ffabffabffabffab;
mem[6851] = 80'h0010ffabffabffabffab;
mem[6852] = 80'h0010ffabffabffabffab;
mem[6853] = 80'h0010ffabffabffabffab;
mem[6854] = 80'h0010ffabffabffabffab;
mem[6855] = 80'h0010ffabffabffabffab;
mem[6856] = 80'h0010ffabffabffabffab;
mem[6857] = 80'h0010ffabffabffabffab;
mem[6858] = 80'h0010ffabffabffabffab;
mem[6859] = 80'h0010ffabffabffabffab;
mem[6860] = 80'h0010ffabffabffabffab;
mem[6861] = 80'h0010ffabffabffabffab;
mem[6862] = 80'h0010ffabffabffabffab;
mem[6863] = 80'h0010ffabffabffabffab;
mem[6864] = 80'h0010ffabffabffabffab;
mem[6865] = 80'h0010ffabffabffabffab;
mem[6866] = 80'h0010ffabffabffabffab;
mem[6867] = 80'h0010ffabffabffabffab;
mem[6868] = 80'h0010ffabffabffabffab;
mem[6869] = 80'h0010ffabffabffabffab;
mem[6870] = 80'h0010ffabffabffabffab;
mem[6871] = 80'h0010ffabffabffabffab;
mem[6872] = 80'h0010ffabffabffabffab;
mem[6873] = 80'h0010ffabffabffabffab;
mem[6874] = 80'h0010ffabffabffabffab;
mem[6875] = 80'h0010ffabffabffabffab;
mem[6876] = 80'h0010ffabffabffabffab;
mem[6877] = 80'h0010ffabffabffabffab;
mem[6878] = 80'h0010ffabffabffabffab;
mem[6879] = 80'h0010ffabffabffabffab;
mem[6880] = 80'h0010ffabffabffabffab;
mem[6881] = 80'h0010ffabffabffabffab;
mem[6882] = 80'h0010ffabffabffabffab;
mem[6883] = 80'h0010ffabffabffabffab;
mem[6884] = 80'h0010ffabffabffabffab;
mem[6885] = 80'h0010ffabffabffabffab;
mem[6886] = 80'h0010ffabffabffabffab;
mem[6887] = 80'h0010ffabffabffabffab;
mem[6888] = 80'h0010ffabffabffabffab;
mem[6889] = 80'h0010ffabffabffabffab;
mem[6890] = 80'h0010ffabffabffabffab;
mem[6891] = 80'h0010ffabffabffabffab;
mem[6892] = 80'h0010ffabffabffabffab;
mem[6893] = 80'h0010ffabffabffabffab;
mem[6894] = 80'h0010ffabffabffabffab;
mem[6895] = 80'h0010ffabffabffabffab;
mem[6896] = 80'h0010ffabffabffabffab;
mem[6897] = 80'h0010ffabffabffabffab;
mem[6898] = 80'h0010ffabffabffabffab;
mem[6899] = 80'h0010ffabffabffabffab;
mem[6900] = 80'h0010ffabffabffabffab;
mem[6901] = 80'h0010ffabffabffabffab;
mem[6902] = 80'h0010ffabffabffabffab;
mem[6903] = 80'h0010ffabffabffabffab;
mem[6904] = 80'h0010ffabffabffabffab;
mem[6905] = 80'h0010ffabffabffabffab;
mem[6906] = 80'h0010ffabffabffabffab;
mem[6907] = 80'h0010ffabffabffabffab;
mem[6908] = 80'h0010ffabffabffabffab;
mem[6909] = 80'h0010ffabffabffabffab;
mem[6910] = 80'h0010ffabffabffabffab;
mem[6911] = 80'h0010ffabffabffabffab;
mem[6912] = 80'h0010ffabffabffabffab;
mem[6913] = 80'h0010ffabffabffabffab;
mem[6914] = 80'h0010ffabffabffabffab;
mem[6915] = 80'h0010ffabffabffabffab;
mem[6916] = 80'h0010ffabffabffabffab;
mem[6917] = 80'h0010ffabffabffabffab;
mem[6918] = 80'h0010ffabffabffabffab;
mem[6919] = 80'h0010ffabffabffabffab;
mem[6920] = 80'h0010ffabffabffabffab;
mem[6921] = 80'h0010ffabffabffabffab;
mem[6922] = 80'h0010ffabffabffabffab;
mem[6923] = 80'h0010ffabffabffabffab;
mem[6924] = 80'h0010ffabffabffabffab;
mem[6925] = 80'h0010ffabffabffabffab;
mem[6926] = 80'h0010ffabffabffabffab;
mem[6927] = 80'h0010ffabffabffabffab;
mem[6928] = 80'h0010ffabffabffabffab;
mem[6929] = 80'h0010ffabffabffabffab;
mem[6930] = 80'h0010ffabffabffabffab;
mem[6931] = 80'h0010ffabffabffabffab;
mem[6932] = 80'h0010ffabffabffabffab;
mem[6933] = 80'h0010ffabffabffabffab;
mem[6934] = 80'h0010ffabffabffabffab;
mem[6935] = 80'h0010ffabffabffabffab;
mem[6936] = 80'h0010ffabffabffabffab;
mem[6937] = 80'h0010ffabffabffabffab;
mem[6938] = 80'h0010ffab2103936275e1;
mem[6939] = 80'h00100231b7d5a94eda40;
mem[6940] = 80'h001072c7a45181094e1d;
mem[6941] = 80'h0112a7fe000000000000;
mem[6942] = 80'h10100000010000010010;
mem[6943] = 80'h00109400000208004500;
mem[6944] = 80'h0010021789df0000fffd;
mem[6945] = 80'h0010adb1c0550102c000;
mem[6946] = 80'h00100001ffabffabffab;
mem[6947] = 80'h0010ffabffabffabffab;
mem[6948] = 80'h0010ffabffabffabffab;
mem[6949] = 80'h0010ffabffabffabffab;
mem[6950] = 80'h0010ffabffabffabffab;
mem[6951] = 80'h0010ffabffabffabffab;
mem[6952] = 80'h0010ffabffabffabffab;
mem[6953] = 80'h0010ffabffabffabffab;
mem[6954] = 80'h0010ffabffabffabffab;
mem[6955] = 80'h0010ffabffabffabffab;
mem[6956] = 80'h0010ffabffabffabffab;
mem[6957] = 80'h0010ffabffabffabffab;
mem[6958] = 80'h0010ffabffabffabffab;
mem[6959] = 80'h0010ffabffabffabffab;
mem[6960] = 80'h0010ffabffabffabffab;
mem[6961] = 80'h0010ffabffabffabffab;
mem[6962] = 80'h0010ffabffabffabffab;
mem[6963] = 80'h0010ffabffabffabffab;
mem[6964] = 80'h0010ffabffabffabffab;
mem[6965] = 80'h0010ffabffabffabffab;
mem[6966] = 80'h0010ffabffabffabffab;
mem[6967] = 80'h0010ffabffabffabffab;
mem[6968] = 80'h0010ffabffabffabffab;
mem[6969] = 80'h0010ffabffabffabffab;
mem[6970] = 80'h0010ffabffabffabffab;
mem[6971] = 80'h0010ffabffabffabffab;
mem[6972] = 80'h0010ffabffabffabffab;
mem[6973] = 80'h0010ffabffabffabffab;
mem[6974] = 80'h0010ffabffabffabffab;
mem[6975] = 80'h0010ffabffabffabffab;
mem[6976] = 80'h0010ffabffabffabffab;
mem[6977] = 80'h0010ffabffabffabffab;
mem[6978] = 80'h0010ffabffabffabffab;
mem[6979] = 80'h0010ffabffabffabffab;
mem[6980] = 80'h0010ffabffabffabffab;
mem[6981] = 80'h0010ffabffabffabffab;
mem[6982] = 80'h0010ffabffabffabffab;
mem[6983] = 80'h0010ffabffabffabffab;
mem[6984] = 80'h0010ffabffabffabffab;
mem[6985] = 80'h0010ffabffabffabffab;
mem[6986] = 80'h0010ffabffabffabffab;
mem[6987] = 80'h0010ffabffabffabffab;
mem[6988] = 80'h0010ffabffabffabffab;
mem[6989] = 80'h0010ffabffabffabffab;
mem[6990] = 80'h0010ffabffabffabffab;
mem[6991] = 80'h0010ffabffabffabffab;
mem[6992] = 80'h0010ffabffabffabffab;
mem[6993] = 80'h0010ffabffabffabffab;
mem[6994] = 80'h0010ffabffabffabffab;
mem[6995] = 80'h0010ffabffabffabffab;
mem[6996] = 80'h0010ffabffabffabffab;
mem[6997] = 80'h0010ffabffabffabffab;
mem[6998] = 80'h0010ffabffabffabffab;
mem[6999] = 80'h0010ffabffabffabffab;
mem[7000] = 80'h0010ffabffabffabffab;
mem[7001] = 80'h0010ffabffabffabffab;
mem[7002] = 80'h0010ffabffabffabffab;
mem[7003] = 80'h0010ffabffabffabffab;
mem[7004] = 80'h0010ffabffabffabffab;
mem[7005] = 80'h0010ffabffabffabffab;
mem[7006] = 80'h0010ffabffabffabffab;
mem[7007] = 80'h0010ffabffabffabffab;
mem[7008] = 80'h0010ff20724d4ead98c0;
mem[7009] = 80'h00108e7c072ea32f9142;
mem[7010] = 80'h001096e73e200712a7f7;
mem[7011] = 80'h01118e00000000000000;
mem[7012] = 80'h10100000010000010010;
mem[7013] = 80'h00109400000208004500;
mem[7014] = 80'h001003fb89e00000fffd;
mem[7015] = 80'h0010abccc0550102c000;
mem[7016] = 80'h00100001ffabffabffab;
mem[7017] = 80'h0010ffabffabffabffab;
mem[7018] = 80'h0010ffabffabffabffab;
mem[7019] = 80'h0010ffabffabffabffab;
mem[7020] = 80'h0010ffabffabffabffab;
mem[7021] = 80'h0010ffabffabffabffab;
mem[7022] = 80'h0010ffabffabffabffab;
mem[7023] = 80'h0010ffabffabffabffab;
mem[7024] = 80'h0010ffabffabffabffab;
mem[7025] = 80'h0010ffabffabffabffab;
mem[7026] = 80'h0010ffabffabffabffab;
mem[7027] = 80'h0010ffabffabffabffab;
mem[7028] = 80'h0010ffabffabffabffab;
mem[7029] = 80'h0010ffabffabffabffab;
mem[7030] = 80'h0010ffabffabffabffab;
mem[7031] = 80'h0010ffabffabffabffab;
mem[7032] = 80'h0010ffabffabffabffab;
mem[7033] = 80'h0010ffabffabffabffab;
mem[7034] = 80'h0010ffabffabffabffab;
mem[7035] = 80'h0010ffabffabffabffab;
mem[7036] = 80'h0010ffabffabffabffab;
mem[7037] = 80'h0010ffabffabffabffab;
mem[7038] = 80'h0010ffabffabffabffab;
mem[7039] = 80'h0010ffabffabffabffab;
mem[7040] = 80'h0010ffabffabffabffab;
mem[7041] = 80'h0010ffabffabffabffab;
mem[7042] = 80'h0010ffabffabffabffab;
mem[7043] = 80'h0010ffabffabffabffab;
mem[7044] = 80'h0010ffabffabffabffab;
mem[7045] = 80'h0010ffabffabffabffab;
mem[7046] = 80'h0010ffabffabffabffab;
mem[7047] = 80'h0010ffabffabffabffab;
mem[7048] = 80'h0010ffabffabffabffab;
mem[7049] = 80'h0010ffabffabffabffab;
mem[7050] = 80'h0010ffabffabffabffab;
mem[7051] = 80'h0010ffabffabffabffab;
mem[7052] = 80'h0010ffabffabffabffab;
mem[7053] = 80'h0010ffabffabffabffab;
mem[7054] = 80'h0010ffabffabffabffab;
mem[7055] = 80'h0010ffabffabffabffab;
mem[7056] = 80'h0010ffabffabffabffab;
mem[7057] = 80'h0010ffabffabffabffab;
mem[7058] = 80'h0010ffabffabffabffab;
mem[7059] = 80'h0010ffabffabffabffab;
mem[7060] = 80'h0010ffabffabffabffab;
mem[7061] = 80'h0010ffabffabffabffab;
mem[7062] = 80'h0010ffabffabffabffab;
mem[7063] = 80'h0010ffabffabffabffab;
mem[7064] = 80'h0010ffabffabffabffab;
mem[7065] = 80'h0010ffabffabffabffab;
mem[7066] = 80'h0010ffabffabffabffab;
mem[7067] = 80'h0010ffabffabffabffab;
mem[7068] = 80'h0010ffabffabffabffab;
mem[7069] = 80'h0010ffabffabffabffab;
mem[7070] = 80'h0010ffabffabffabffab;
mem[7071] = 80'h0010ffabffabffabffab;
mem[7072] = 80'h0010ffabffabffabffab;
mem[7073] = 80'h0010ffabffabffabffab;
mem[7074] = 80'h0010ffabffabffabffab;
mem[7075] = 80'h0010ffabffabffabffab;
mem[7076] = 80'h0010ffabffabffabffab;
mem[7077] = 80'h0010ffabffabffabffab;
mem[7078] = 80'h0010ffabffabffabffab;
mem[7079] = 80'h0010ffabffabffabffab;
mem[7080] = 80'h0010ffabffabffabffab;
mem[7081] = 80'h0010ffabffabffabffab;
mem[7082] = 80'h0010ffabffabffabffab;
mem[7083] = 80'h0010ffabffabffabffab;
mem[7084] = 80'h0010ffabffabffabffab;
mem[7085] = 80'h0010ffabffabffabffab;
mem[7086] = 80'h0010ffabffabffabffab;
mem[7087] = 80'h0010ffabffabffabffab;
mem[7088] = 80'h0010ffabffabffabffab;
mem[7089] = 80'h0010ffabffabffabffab;
mem[7090] = 80'h0010ffabffabffabffab;
mem[7091] = 80'h0010ffabffabffabffab;
mem[7092] = 80'h0010ffabffabffabffab;
mem[7093] = 80'h0010ffabffabffabffab;
mem[7094] = 80'h0010ffabffabffabffab;
mem[7095] = 80'h0010ffabffabffabffab;
mem[7096] = 80'h0010ffabffabffabffab;
mem[7097] = 80'h0010ffabffabffabffab;
mem[7098] = 80'h0010ffabffabffabffab;
mem[7099] = 80'h0010ffabffabffabffab;
mem[7100] = 80'h0010ffabffabffabffab;
mem[7101] = 80'h0010ffabffabffabffab;
mem[7102] = 80'h0010ffabffabffabffab;
mem[7103] = 80'h0010ffabffabffabffab;
mem[7104] = 80'h0010ffabffabffabffab;
mem[7105] = 80'h0010ffabffabffabffab;
mem[7106] = 80'h0010ffabffabffabffab;
mem[7107] = 80'h0010ffabffabffabffab;
mem[7108] = 80'h0010ffabffabffabffab;
mem[7109] = 80'h0010ffabffabffabffab;
mem[7110] = 80'h0010ffabffabffabffab;
mem[7111] = 80'h0010ffabffabffabffab;
mem[7112] = 80'h0010ffabffabffabffab;
mem[7113] = 80'h0010ffabffabffabffab;
mem[7114] = 80'h0010ffabffabffabffab;
mem[7115] = 80'h0010ffabffabffabffab;
mem[7116] = 80'h0010ffabffabffabffab;
mem[7117] = 80'h0010ffabffabffabffab;
mem[7118] = 80'h0010ffabffabffabffab;
mem[7119] = 80'h0010ffabffabffabffab;
mem[7120] = 80'h0010ffabffabffabffab;
mem[7121] = 80'h0010ffabffabffabffab;
mem[7122] = 80'h0010ffabffabffabffab;
mem[7123] = 80'h0010ffabffabffabffab;
mem[7124] = 80'h0010ffabffabffabffab;
mem[7125] = 80'h0010ffabffabffabffab;
mem[7126] = 80'h0010ffabffabffabffab;
mem[7127] = 80'h0010ffabffabffabffab;
mem[7128] = 80'h0010ffabffabffabffab;
mem[7129] = 80'h0010ffabffabffabffab;
mem[7130] = 80'h0010ffabffabffabffab;
mem[7131] = 80'h0010ffabffabffabffab;
mem[7132] = 80'h0010ffabffabffabffab;
mem[7133] = 80'h0010ffabffabffabffab;
mem[7134] = 80'h0010ffabffabffabffab;
mem[7135] = 80'h0010ffabffabffabffab;
mem[7136] = 80'h0010ffabffabffabffab;
mem[7137] = 80'h0010ffabffabffabffab;
mem[7138] = 80'h0010ffabffabff1f0170;
mem[7139] = 80'h0010de2c51f1b4c84232;
mem[7140] = 80'h0010430195df0d9c82da;
mem[7141] = 80'h01156e32e13b82000000;
mem[7142] = 80'h10100000010000010010;
mem[7143] = 80'h00109400000208004500;
mem[7144] = 80'h0010021689e10000fffd;
mem[7145] = 80'h0010adb0c0550102c000;
mem[7146] = 80'h00100001ffabffabffab;
mem[7147] = 80'h0010ffabffabffabffab;
mem[7148] = 80'h0010ffabffabffabffab;
mem[7149] = 80'h0010ffabffabffabffab;
mem[7150] = 80'h0010ffabffabffabffab;
mem[7151] = 80'h0010ffabffabffabffab;
mem[7152] = 80'h0010ffabffabffabffab;
mem[7153] = 80'h0010ffabffabffabffab;
mem[7154] = 80'h0010ffabffabffabffab;
mem[7155] = 80'h0010ffabffabffabffab;
mem[7156] = 80'h0010ffabffabffabffab;
mem[7157] = 80'h0010ffabffabffabffab;
mem[7158] = 80'h0010ffabffabffabffab;
mem[7159] = 80'h0010ffabffabffabffab;
mem[7160] = 80'h0010ffabffabffabffab;
mem[7161] = 80'h0010ffabffabffabffab;
mem[7162] = 80'h0010ffabffabffabffab;
mem[7163] = 80'h0010ffabffabffabffab;
mem[7164] = 80'h0010ffabffabffabffab;
mem[7165] = 80'h0010ffabffabffabffab;
mem[7166] = 80'h0010ffabffabffabffab;
mem[7167] = 80'h0010ffabffabffabffab;
mem[7168] = 80'h0010ffabffabffabffab;
mem[7169] = 80'h0010ffabffabffabffab;
mem[7170] = 80'h0010ffabffabffabffab;
mem[7171] = 80'h0010ffabffabffabffab;
mem[7172] = 80'h0010ffabffabffabffab;
mem[7173] = 80'h0010ffabffabffabffab;
mem[7174] = 80'h0010ffabffabffabffab;
mem[7175] = 80'h0010ffabffabffabffab;
mem[7176] = 80'h0010ffabffabffabffab;
mem[7177] = 80'h0010ffabffabffabffab;
mem[7178] = 80'h0010ffabffabffabffab;
mem[7179] = 80'h0010ffabffabffabffab;
mem[7180] = 80'h0010ffabffabffabffab;
mem[7181] = 80'h0010ffabffabffabffab;
mem[7182] = 80'h0010ffabffabffabffab;
mem[7183] = 80'h0010ffabffabffabffab;
mem[7184] = 80'h0010ffabffabffabffab;
mem[7185] = 80'h0010ffabffabffabffab;
mem[7186] = 80'h0010ffabffabffabffab;
mem[7187] = 80'h0010ffabffabffabffab;
mem[7188] = 80'h0010ffabffabffabffab;
mem[7189] = 80'h0010ffabffabffabffab;
mem[7190] = 80'h0010ffabffabffabffab;
mem[7191] = 80'h0010ffabffabffabffab;
mem[7192] = 80'h0010ffabffabffabffab;
mem[7193] = 80'h0010ffabffabffabffab;
mem[7194] = 80'h0010ffabffabffabffab;
mem[7195] = 80'h0010ffabffabffabffab;
mem[7196] = 80'h0010ffabffabffabffab;
mem[7197] = 80'h0010ffabffabffabffab;
mem[7198] = 80'h0010ffabffabffabffab;
mem[7199] = 80'h0010ffabffabffabffab;
mem[7200] = 80'h0010ffabffabffabffab;
mem[7201] = 80'h0010ffabffabffabffab;
mem[7202] = 80'h0010ffabffabffabffab;
mem[7203] = 80'h0010ffabffabffabffab;
mem[7204] = 80'h0010ffabffabffabffab;
mem[7205] = 80'h0010ffabffabffabffab;
mem[7206] = 80'h0010ffabffabffabffab;
mem[7207] = 80'h0010ffabffabffabffab;
mem[7208] = 80'h00101e70aef2f428330b;
mem[7209] = 80'h00100390b5aef444d65c;
mem[7210] = 80'h011060e026a8b7f1750c;
mem[7211] = 80'h10100000010000010010;
mem[7212] = 80'h00109400000208004500;
mem[7213] = 80'h001003f989e20000fffd;
mem[7214] = 80'h0010abccc0550102c000;
mem[7215] = 80'h00100001ffabffabffab;
mem[7216] = 80'h0010ffabffabffabffab;
mem[7217] = 80'h0010ffabffabffabffab;
mem[7218] = 80'h0010ffabffabffabffab;
mem[7219] = 80'h0010ffabffabffabffab;
mem[7220] = 80'h0010ffabffabffabffab;
mem[7221] = 80'h0010ffabffabffabffab;
mem[7222] = 80'h0010ffabffabffabffab;
mem[7223] = 80'h0010ffabffabffabffab;
mem[7224] = 80'h0010ffabffabffabffab;
mem[7225] = 80'h0010ffabffabffabffab;
mem[7226] = 80'h0010ffabffabffabffab;
mem[7227] = 80'h0010ffabffabffabffab;
mem[7228] = 80'h0010ffabffabffabffab;
mem[7229] = 80'h0010ffabffabffabffab;
mem[7230] = 80'h0010ffabffabffabffab;
mem[7231] = 80'h0010ffabffabffabffab;
mem[7232] = 80'h0010ffabffabffabffab;
mem[7233] = 80'h0010ffabffabffabffab;
mem[7234] = 80'h0010ffabffabffabffab;
mem[7235] = 80'h0010ffabffabffabffab;
mem[7236] = 80'h0010ffabffabffabffab;
mem[7237] = 80'h0010ffabffabffabffab;
mem[7238] = 80'h0010ffabffabffabffab;
mem[7239] = 80'h0010ffabffabffabffab;
mem[7240] = 80'h0010ffabffabffabffab;
mem[7241] = 80'h0010ffabffabffabffab;
mem[7242] = 80'h0010ffabffabffabffab;
mem[7243] = 80'h0010ffabffabffabffab;
mem[7244] = 80'h0010ffabffabffabffab;
mem[7245] = 80'h0010ffabffabffabffab;
mem[7246] = 80'h0010ffabffabffabffab;
mem[7247] = 80'h0010ffabffabffabffab;
mem[7248] = 80'h0010ffabffabffabffab;
mem[7249] = 80'h0010ffabffabffabffab;
mem[7250] = 80'h0010ffabffabffabffab;
mem[7251] = 80'h0010ffabffabffabffab;
mem[7252] = 80'h0010ffabffabffabffab;
mem[7253] = 80'h0010ffabffabffabffab;
mem[7254] = 80'h0010ffabffabffabffab;
mem[7255] = 80'h0010ffabffabffabffab;
mem[7256] = 80'h0010ffabffabffabffab;
mem[7257] = 80'h0010ffabffabffabffab;
mem[7258] = 80'h0010ffabffabffabffab;
mem[7259] = 80'h0010ffabffabffabffab;
mem[7260] = 80'h0010ffabffabffabffab;
mem[7261] = 80'h0010ffabffabffabffab;
mem[7262] = 80'h0010ffabffabffabffab;
mem[7263] = 80'h0010ffabffabffabffab;
mem[7264] = 80'h0010ffabffabffabffab;
mem[7265] = 80'h0010ffabffabffabffab;
mem[7266] = 80'h0010ffabffabffabffab;
mem[7267] = 80'h0010ffabffabffabffab;
mem[7268] = 80'h0010ffabffabffabffab;
mem[7269] = 80'h0010ffabffabffabffab;
mem[7270] = 80'h0010ffabffabffabffab;
mem[7271] = 80'h0010ffabffabffabffab;
mem[7272] = 80'h0010ffabffabffabffab;
mem[7273] = 80'h0010ffabffabffabffab;
mem[7274] = 80'h0010ffabffabffabffab;
mem[7275] = 80'h0010ffabffabffabffab;
mem[7276] = 80'h0010ffabffabffabffab;
mem[7277] = 80'h0010ffabffabffabffab;
mem[7278] = 80'h0010ffabffabffabffab;
mem[7279] = 80'h0010ffabffabffabffab;
mem[7280] = 80'h0010ffabffabffabffab;
mem[7281] = 80'h0010ffabffabffabffab;
mem[7282] = 80'h0010ffabffabffabffab;
mem[7283] = 80'h0010ffabffabffabffab;
mem[7284] = 80'h0010ffabffabffabffab;
mem[7285] = 80'h0010ffabffabffabffab;
mem[7286] = 80'h0010ffabffabffabffab;
mem[7287] = 80'h0010ffabffabffabffab;
mem[7288] = 80'h0010ffabffabffabffab;
mem[7289] = 80'h0010ffabffabffabffab;
mem[7290] = 80'h0010ffabffabffabffab;
mem[7291] = 80'h0010ffabffabffabffab;
mem[7292] = 80'h0010ffabffabffabffab;
mem[7293] = 80'h0010ffabffabffabffab;
mem[7294] = 80'h0010ffabffabffabffab;
mem[7295] = 80'h0010ffabffabffabffab;
mem[7296] = 80'h0010ffabffabffabffab;
mem[7297] = 80'h0010ffabffabffabffab;
mem[7298] = 80'h0010ffabffabffabffab;
mem[7299] = 80'h0010ffabffabffabffab;
mem[7300] = 80'h0010ffabffabffabffab;
mem[7301] = 80'h0010ffabffabffabffab;
mem[7302] = 80'h0010ffabffabffabffab;
mem[7303] = 80'h0010ffabffabffabffab;
mem[7304] = 80'h0010ffabffabffabffab;
mem[7305] = 80'h0010ffabffabffabffab;
mem[7306] = 80'h0010ffabffabffabffab;
mem[7307] = 80'h0010ffabffabffabffab;
mem[7308] = 80'h0010ffabffabffabffab;
mem[7309] = 80'h0010ffabffabffabffab;
mem[7310] = 80'h0010ffabffabffabffab;
mem[7311] = 80'h0010ffabffabffabffab;
mem[7312] = 80'h0010ffabffabffabffab;
mem[7313] = 80'h0010ffabffabffabffab;
mem[7314] = 80'h0010ffabffabffabffab;
mem[7315] = 80'h0010ffabffabffabffab;
mem[7316] = 80'h0010ffabffabffabffab;
mem[7317] = 80'h0010ffabffabffabffab;
mem[7318] = 80'h0010ffabffabffabffab;
mem[7319] = 80'h0010ffabffabffabffab;
mem[7320] = 80'h0010ffabffabffabffab;
mem[7321] = 80'h0010ffabffabffabffab;
mem[7322] = 80'h0010ffabffabffabffab;
mem[7323] = 80'h0010ffabffabffabffab;
mem[7324] = 80'h0010ffabffabffabffab;
mem[7325] = 80'h0010ffabffabffabffab;
mem[7326] = 80'h0010ffabffabffabffab;
mem[7327] = 80'h0010ffabffabffabffab;
mem[7328] = 80'h0010ffabffabffabffab;
mem[7329] = 80'h0010ffabffabffabffab;
mem[7330] = 80'h0010ffabffabffabffab;
mem[7331] = 80'h0010ffabffabffabffab;
mem[7332] = 80'h0010ffabffabffabffab;
mem[7333] = 80'h0010ffabffabffabffab;
mem[7334] = 80'h0010ffabffabffabffab;
mem[7335] = 80'h0010ffabffabffabffab;
mem[7336] = 80'h0010ffabffabffabffab;
mem[7337] = 80'h0010ffabff1de2cc879c;
mem[7338] = 80'h0010a274cb5fe73d98ea;
mem[7339] = 80'h00103701ae377f4343bc;
mem[7340] = 80'h0113a1c6e30000000000;
mem[7341] = 80'h10100000010000010010;
mem[7342] = 80'h00109400000208004500;
mem[7343] = 80'h0010021389e30000fffd;
mem[7344] = 80'h0010adb1c0550102c000;
mem[7345] = 80'h00100001ffabffabffab;
mem[7346] = 80'h0010ffabffabffabffab;
mem[7347] = 80'h0010ffabffabffabffab;
mem[7348] = 80'h0010ffabffabffabffab;
mem[7349] = 80'h0010ffabffabffabffab;
mem[7350] = 80'h0010ffabffabffabffab;
mem[7351] = 80'h0010ffabffabffabffab;
mem[7352] = 80'h0010ffabffabffabffab;
mem[7353] = 80'h0010ffabffabffabffab;
mem[7354] = 80'h0010ffabffabffabffab;
mem[7355] = 80'h0010ffabffabffabffab;
mem[7356] = 80'h0010ffabffabffabffab;
mem[7357] = 80'h0010ffabffabffabffab;
mem[7358] = 80'h0010ffabffabffabffab;
mem[7359] = 80'h0010ffabffabffabffab;
mem[7360] = 80'h0010ffabffabffabffab;
mem[7361] = 80'h0010ffabffabffabffab;
mem[7362] = 80'h0010ffabffabffabffab;
mem[7363] = 80'h0010ffabffabffabffab;
mem[7364] = 80'h0010ffabffabffabffab;
mem[7365] = 80'h0010ffabffabffabffab;
mem[7366] = 80'h0010ffabffabffabffab;
mem[7367] = 80'h0010ffabffabffabffab;
mem[7368] = 80'h0010ffabffabffabffab;
mem[7369] = 80'h0010ffabffabffabffab;
mem[7370] = 80'h0010ffabffabffabffab;
mem[7371] = 80'h0010ffabffabffabffab;
mem[7372] = 80'h0010ffabffabffabffab;
mem[7373] = 80'h0010ffabffabffabffab;
mem[7374] = 80'h0010ffabffabffabffab;
mem[7375] = 80'h0010ffabffabffabffab;
mem[7376] = 80'h0010ffabffabffabffab;
mem[7377] = 80'h0010ffabffabffabffab;
mem[7378] = 80'h0010ffabffabffabffab;
mem[7379] = 80'h0010ffabffabffabffab;
mem[7380] = 80'h0010ffabffabffabffab;
mem[7381] = 80'h0010ffabffabffabffab;
mem[7382] = 80'h0010ffabffabffabffab;
mem[7383] = 80'h0010ffabffabffabffab;
mem[7384] = 80'h0010ffabffabffabffab;
mem[7385] = 80'h0010ffabffabffabffab;
mem[7386] = 80'h0010ffabffabffabffab;
mem[7387] = 80'h0010ffabffabffabffab;
mem[7388] = 80'h0010ffabffabffabffab;
mem[7389] = 80'h0010ffabffabffabffab;
mem[7390] = 80'h0010ffabffabffabffab;
mem[7391] = 80'h0010ffabffabffabffab;
mem[7392] = 80'h0010ffabffabffabffab;
mem[7393] = 80'h0010ffabffabffabffab;
mem[7394] = 80'h0010ffabffabffabffab;
mem[7395] = 80'h0010ffabffabffabffab;
mem[7396] = 80'h0010ffabffabffabffab;
mem[7397] = 80'h0010ffabffabffabffab;
mem[7398] = 80'h0010ffabffabffabffab;
mem[7399] = 80'h0010ffabffabffabffab;
mem[7400] = 80'h0010ffabffabffabffab;
mem[7401] = 80'h0010ffabffabffabffab;
mem[7402] = 80'h0010ffabffabffabffab;
mem[7403] = 80'h0010ffabffabffabffab;
mem[7404] = 80'h0010ffabffabffabffab;
mem[7405] = 80'h0010ffabffabffabffab;
mem[7406] = 80'h0010ffabffabff1c9312;
mem[7407] = 80'h0010ab44dbb6749435ba;
mem[7408] = 80'h0010751fe612ff27a52c;
mem[7409] = 80'h01153c987e9b03000000;
mem[7410] = 80'h10100000010000010010;
mem[7411] = 80'h00109400000208004500;
mem[7412] = 80'h001003f989e40000fffd;
mem[7413] = 80'h0010abcac0550102c000;
mem[7414] = 80'h00100001ffabffabffab;
mem[7415] = 80'h0010ffabffabffabffab;
mem[7416] = 80'h0010ffabffabffabffab;
mem[7417] = 80'h0010ffabffabffabffab;
mem[7418] = 80'h0010ffabffabffabffab;
mem[7419] = 80'h0010ffabffabffabffab;
mem[7420] = 80'h0010ffabffabffabffab;
mem[7421] = 80'h0010ffabffabffabffab;
mem[7422] = 80'h0010ffabffabffabffab;
mem[7423] = 80'h0010ffabffabffabffab;
mem[7424] = 80'h0010ffabffabffabffab;
mem[7425] = 80'h0010ffabffabffabffab;
mem[7426] = 80'h0010ffabffabffabffab;
mem[7427] = 80'h0010ffabffabffabffab;
mem[7428] = 80'h0010ffabffabffabffab;
mem[7429] = 80'h0010ffabffabffabffab;
mem[7430] = 80'h0010ffabffabffabffab;
mem[7431] = 80'h0010ffabffabffabffab;
mem[7432] = 80'h0010ffabffabffabffab;
mem[7433] = 80'h0010ffabffabffabffab;
mem[7434] = 80'h0010ffabffabffabffab;
mem[7435] = 80'h0010ffabffabffabffab;
mem[7436] = 80'h0010ffabffabffabffab;
mem[7437] = 80'h0010ffabffabffabffab;
mem[7438] = 80'h0010ffabffabffabffab;
mem[7439] = 80'h0010ffabffabffabffab;
mem[7440] = 80'h0010ffabffabffabffab;
mem[7441] = 80'h0010ffabffabffabffab;
mem[7442] = 80'h0010ffabffabffabffab;
mem[7443] = 80'h0010ffabffabffabffab;
mem[7444] = 80'h0010ffabffabffabffab;
mem[7445] = 80'h0010ffabffabffabffab;
mem[7446] = 80'h0010ffabffabffabffab;
mem[7447] = 80'h0010ffabffabffabffab;
mem[7448] = 80'h0010ffabffabffabffab;
mem[7449] = 80'h0010ffabffabffabffab;
mem[7450] = 80'h0010ffabffabffabffab;
mem[7451] = 80'h0010ffabffabffabffab;
mem[7452] = 80'h0010ffabffabffabffab;
mem[7453] = 80'h0010ffabffabffabffab;
mem[7454] = 80'h0010ffabffabffabffab;
mem[7455] = 80'h0010ffabffabffabffab;
mem[7456] = 80'h0010ffabffabffabffab;
mem[7457] = 80'h0010ffabffabffabffab;
mem[7458] = 80'h0010ffabffabffabffab;
mem[7459] = 80'h0010ffabffabffabffab;
mem[7460] = 80'h0010ffabffabffabffab;
mem[7461] = 80'h0010ffabffabffabffab;
mem[7462] = 80'h0010ffabffabffabffab;
mem[7463] = 80'h0010ffabffabffabffab;
mem[7464] = 80'h0010ffabffabffabffab;
mem[7465] = 80'h0010ffabffabffabffab;
mem[7466] = 80'h0010ffabffabffabffab;
mem[7467] = 80'h0010ffabffabffabffab;
mem[7468] = 80'h0010ffabffabffabffab;
mem[7469] = 80'h0010ffabffabffabffab;
mem[7470] = 80'h0010ffabffabffabffab;
mem[7471] = 80'h0010ffabffabffabffab;
mem[7472] = 80'h0010ffabffabffabffab;
mem[7473] = 80'h0010ffabffabffabffab;
mem[7474] = 80'h0010ffabffabffabffab;
mem[7475] = 80'h0010ffabffabffabffab;
mem[7476] = 80'h0010ffabffabffabffab;
mem[7477] = 80'h0010ffabffabffabffab;
mem[7478] = 80'h0010ffabffabffabffab;
mem[7479] = 80'h0010ffabffabffabffab;
mem[7480] = 80'h0010ffabffabffabffab;
mem[7481] = 80'h0010ffabffabffabffab;
mem[7482] = 80'h0010ffabffabffabffab;
mem[7483] = 80'h0010ffabffabffabffab;
mem[7484] = 80'h0010ffabffabffabffab;
mem[7485] = 80'h0010ffabffabffabffab;
mem[7486] = 80'h0010ffabffabffabffab;
mem[7487] = 80'h0010ffabffabffabffab;
mem[7488] = 80'h0010ffabffabffabffab;
mem[7489] = 80'h0010ffabffabffabffab;
mem[7490] = 80'h0010ffabffabffabffab;
mem[7491] = 80'h0010ffabffabffabffab;
mem[7492] = 80'h0010ffabffabffabffab;
mem[7493] = 80'h0010ffabffabffabffab;
mem[7494] = 80'h0010ffabffabffabffab;
mem[7495] = 80'h0010ffabffabffabffab;
mem[7496] = 80'h0010ffabffabffabffab;
mem[7497] = 80'h0010ffabffabffabffab;
mem[7498] = 80'h0010ffabffabffabffab;
mem[7499] = 80'h0010ffabffabffabffab;
mem[7500] = 80'h0010ffabffabffabffab;
mem[7501] = 80'h0010ffabffabffabffab;
mem[7502] = 80'h0010ffabffabffabffab;
mem[7503] = 80'h0010ffabffabffabffab;
mem[7504] = 80'h0010ffabffabffabffab;
mem[7505] = 80'h0010ffabffabffabffab;
mem[7506] = 80'h0010ffabffabffabffab;
mem[7507] = 80'h0010ffabffabffabffab;
mem[7508] = 80'h0010ffabffabffabffab;
mem[7509] = 80'h0010ffabffabffabffab;
mem[7510] = 80'h0010ffabffabffabffab;
mem[7511] = 80'h0010ffabffabffabffab;
mem[7512] = 80'h0010ffabffabffabffab;
mem[7513] = 80'h0010ffabffabffabffab;
mem[7514] = 80'h0010ffabffabffabffab;
mem[7515] = 80'h0010ffabffabffabffab;
mem[7516] = 80'h0010ffabffabffabffab;
mem[7517] = 80'h0010ffabffabffabffab;
mem[7518] = 80'h0010ffabffabffabffab;
mem[7519] = 80'h0010ffabffabffabffab;
mem[7520] = 80'h0010ffabffabffabffab;
mem[7521] = 80'h0010ffabffabffabffab;
mem[7522] = 80'h0010ffabffabffabffab;
mem[7523] = 80'h0010ffabffabffabffab;
mem[7524] = 80'h0010ffabffabffabffab;
mem[7525] = 80'h0010ffabffabffabffab;
mem[7526] = 80'h0010ffabffabffabffab;
mem[7527] = 80'h0010ffabffabffabffab;
mem[7528] = 80'h0010ffabffabffabffab;
mem[7529] = 80'h0010ffabffabffabffab;
mem[7530] = 80'h0010ffabffabffabffab;
mem[7531] = 80'h0010ffabffabffabffab;
mem[7532] = 80'h0010ffabffabffabffab;
mem[7533] = 80'h0010ffabffabffabffab;
mem[7534] = 80'h0010ffabffabffabffab;
mem[7535] = 80'h0010ffabffabffabffab;
mem[7536] = 80'h0010ffabff1bb7d64195;
mem[7537] = 80'h0010cf39f42cdaab1923;
mem[7538] = 80'h001000041a4ebff075d0;
mem[7539] = 80'h011371d58b0000000000;
mem[7540] = 80'h10100000010000010010;
mem[7541] = 80'h00109400000208004500;
mem[7542] = 80'h0010021289e50000fffd;
mem[7543] = 80'h0010adb0c0550102c000;
mem[7544] = 80'h00100001ffabffabffab;
mem[7545] = 80'h0010ffabffabffabffab;
mem[7546] = 80'h0010ffabffabffabffab;
mem[7547] = 80'h0010ffabffabffabffab;
mem[7548] = 80'h0010ffabffabffabffab;
mem[7549] = 80'h0010ffabffabffabffab;
mem[7550] = 80'h0010ffabffabffabffab;
mem[7551] = 80'h0010ffabffabffabffab;
mem[7552] = 80'h0010ffabffabffabffab;
mem[7553] = 80'h0010ffabffabffabffab;
mem[7554] = 80'h0010ffabffabffabffab;
mem[7555] = 80'h0010ffabffabffabffab;
mem[7556] = 80'h0010ffabffabffabffab;
mem[7557] = 80'h0010ffabffabffabffab;
mem[7558] = 80'h0010ffabffabffabffab;
mem[7559] = 80'h0010ffabffabffabffab;
mem[7560] = 80'h0010ffabffabffabffab;
mem[7561] = 80'h0010ffabffabffabffab;
mem[7562] = 80'h0010ffabffabffabffab;
mem[7563] = 80'h0010ffabffabffabffab;
mem[7564] = 80'h0010ffabffabffabffab;
mem[7565] = 80'h0010ffabffabffabffab;
mem[7566] = 80'h0010ffabffabffabffab;
mem[7567] = 80'h0010ffabffabffabffab;
mem[7568] = 80'h0010ffabffabffabffab;
mem[7569] = 80'h0010ffabffabffabffab;
mem[7570] = 80'h0010ffabffabffabffab;
mem[7571] = 80'h0010ffabffabffabffab;
mem[7572] = 80'h0010ffabffabffabffab;
mem[7573] = 80'h0010ffabffabffabffab;
mem[7574] = 80'h0010ffabffabffabffab;
mem[7575] = 80'h0010ffabffabffabffab;
mem[7576] = 80'h0010ffabffabffabffab;
mem[7577] = 80'h0010ffabffabffabffab;
mem[7578] = 80'h0010ffabffabffabffab;
mem[7579] = 80'h0010ffabffabffabffab;
mem[7580] = 80'h0010ffabffabffabffab;
mem[7581] = 80'h0010ffabffabffabffab;
mem[7582] = 80'h0010ffabffabffabffab;
mem[7583] = 80'h0010ffabffabffabffab;
mem[7584] = 80'h0010ffabffabffabffab;
mem[7585] = 80'h0010ffabffabffabffab;
mem[7586] = 80'h0010ffabffabffabffab;
mem[7587] = 80'h0010ffabffabffabffab;
mem[7588] = 80'h0010ffabffabffabffab;
mem[7589] = 80'h0010ffabffabffabffab;
mem[7590] = 80'h0010ffabffabffabffab;
mem[7591] = 80'h0010ffabffabffabffab;
mem[7592] = 80'h0010ffabffabffabffab;
mem[7593] = 80'h0010ffabffabffabffab;
mem[7594] = 80'h0010ffabffabffabffab;
mem[7595] = 80'h0010ffabffabffabffab;
mem[7596] = 80'h0010ffabffabffabffab;
mem[7597] = 80'h0010ffabffabffabffab;
mem[7598] = 80'h0010ffabffabffabffab;
mem[7599] = 80'h0010ffabffabffabffab;
mem[7600] = 80'h0010ffabffabffabffab;
mem[7601] = 80'h0010ffabffabffabffab;
mem[7602] = 80'h0010ffabffabffabffab;
mem[7603] = 80'h0010ffabffabffabffab;
mem[7604] = 80'h0010ffabffabffabffab;
mem[7605] = 80'h0010ffabffab1ac6086d;
mem[7606] = 80'h00104db6fb4be7082cf4;
mem[7607] = 80'h0010d6d1304bc114b79b;
mem[7608] = 80'h0114851b855100000000;
mem[7609] = 80'h10100000010000010010;
mem[7610] = 80'h00109400000208004500;
mem[7611] = 80'h0010012089e60000fffd;
mem[7612] = 80'h0010aea1c0550102c000;
mem[7613] = 80'h00100001ffabffabffab;
mem[7614] = 80'h0010ffabffabffabffab;
mem[7615] = 80'h0010ffabffabffabffab;
mem[7616] = 80'h0010ffabffabffabffab;
mem[7617] = 80'h0010ffabffabffabffab;
mem[7618] = 80'h0010ffabffabffabffab;
mem[7619] = 80'h0010ffabffabffabffab;
mem[7620] = 80'h0010ffabffabffabffab;
mem[7621] = 80'h0010ffabffabffabffab;
mem[7622] = 80'h0010ffabffabffabffab;
mem[7623] = 80'h0010ffabffabffabffab;
mem[7624] = 80'h0010ffabffabffabffab;
mem[7625] = 80'h0010ffabffabffabffab;
mem[7626] = 80'h0010ffabffabffabffab;
mem[7627] = 80'h0010ffabffabffabffab;
mem[7628] = 80'h0010ffabffabffabffab;
mem[7629] = 80'h0010ffabffabffabffab;
mem[7630] = 80'h0010ffabffabffabffab;
mem[7631] = 80'h0010ffabffabffabffab;
mem[7632] = 80'h0010ffabffabffabffab;
mem[7633] = 80'h0010ffabffabffabffab;
mem[7634] = 80'h0010ffabffabffabffab;
mem[7635] = 80'h0010ffabffabffabffab;
mem[7636] = 80'h0010ffabffabffabffab;
mem[7637] = 80'h0010ffabffabffabffab;
mem[7638] = 80'h0010ffabffabffabffab;
mem[7639] = 80'h0010ffabffabffabffab;
mem[7640] = 80'h0010ffabffabffabffab;
mem[7641] = 80'h0010ffabffabffabffab;
mem[7642] = 80'h0010ffabffabffabffab;
mem[7643] = 80'h0010ffabffabffabffab;
mem[7644] = 80'h0010ffab19546a18253c;
mem[7645] = 80'h0010bc8bbb7fa4c2c8a2;
mem[7646] = 80'h0010c1b93acb75611fc3;
mem[7647] = 80'h01125ac1000000000000;
mem[7648] = 80'h10100000010000010010;
mem[7649] = 80'h00109400000208004500;
mem[7650] = 80'h001000a789e70000fffd;
mem[7651] = 80'h0010af19c0550102c000;
mem[7652] = 80'h00100001ffabffabffab;
mem[7653] = 80'h0010ffabffabffabffab;
mem[7654] = 80'h0010ffabffabffabffab;
mem[7655] = 80'h0010ffabffabffabffab;
mem[7656] = 80'h0010ffabffabffabffab;
mem[7657] = 80'h0010ffabffabffabffab;
mem[7658] = 80'h0010ffabffabffabffab;
mem[7659] = 80'h0010ffabffabffabffab;
mem[7660] = 80'h0010ffabffabffabffab;
mem[7661] = 80'h0010ffabffabffabffab;
mem[7662] = 80'h0010ffabffabffabffab;
mem[7663] = 80'h0010ffabffabffabffab;
mem[7664] = 80'h0010ffabffabffabffab;
mem[7665] = 80'h0010ffabffabffabffab;
mem[7666] = 80'h0010ffabffabffabffab;
mem[7667] = 80'h0010ffabffabffabffab;
mem[7668] = 80'h0010ff1825b434fd457e;
mem[7669] = 80'h00103470ad232f3d721b;
mem[7670] = 80'h0010e8b1ed1907f1915b;
mem[7671] = 80'h0111eb00000000000000;
mem[7672] = 80'h10100000010000010010;
mem[7673] = 80'h00109400000208004500;
mem[7674] = 80'h0010034389e80000fffd;
mem[7675] = 80'h0010ac7cc0550102c000;
mem[7676] = 80'h00100001ffabffabffab;
mem[7677] = 80'h0010ffabffabffabffab;
mem[7678] = 80'h0010ffabffabffabffab;
mem[7679] = 80'h0010ffabffabffabffab;
mem[7680] = 80'h0010ffabffabffabffab;
mem[7681] = 80'h0010ffabffabffabffab;
mem[7682] = 80'h0010ffabffabffabffab;
mem[7683] = 80'h0010ffabffabffabffab;
mem[7684] = 80'h0010ffabffabffabffab;
mem[7685] = 80'h0010ffabffabffabffab;
mem[7686] = 80'h0010ffabffabffabffab;
mem[7687] = 80'h0010ffabffabffabffab;
mem[7688] = 80'h0010ffabffabffabffab;
mem[7689] = 80'h0010ffabffabffabffab;
mem[7690] = 80'h0010ffabffabffabffab;
mem[7691] = 80'h0010ffabffabffabffab;
mem[7692] = 80'h0010ffabffabffabffab;
mem[7693] = 80'h0010ffabffabffabffab;
mem[7694] = 80'h0010ffabffabffabffab;
mem[7695] = 80'h0010ffabffabffabffab;
mem[7696] = 80'h0010ffabffabffabffab;
mem[7697] = 80'h0010ffabffabffabffab;
mem[7698] = 80'h0010ffabffabffabffab;
mem[7699] = 80'h0010ffabffabffabffab;
mem[7700] = 80'h0010ffabffabffabffab;
mem[7701] = 80'h0010ffabffabffabffab;
mem[7702] = 80'h0010ffabffabffabffab;
mem[7703] = 80'h0010ffabffabffabffab;
mem[7704] = 80'h0010ffabffabffabffab;
mem[7705] = 80'h0010ffabffabffabffab;
mem[7706] = 80'h0010ffabffabffabffab;
mem[7707] = 80'h0010ffabffabffabffab;
mem[7708] = 80'h0010ffabffabffabffab;
mem[7709] = 80'h0010ffabffabffabffab;
mem[7710] = 80'h0010ffabffabffabffab;
mem[7711] = 80'h0010ffabffabffabffab;
mem[7712] = 80'h0010ffabffabffabffab;
mem[7713] = 80'h0010ffabffabffabffab;
mem[7714] = 80'h0010ffabffabffabffab;
mem[7715] = 80'h0010ffabffabffabffab;
mem[7716] = 80'h0010ffabffabffabffab;
mem[7717] = 80'h0010ffabffabffabffab;
mem[7718] = 80'h0010ffabffabffabffab;
mem[7719] = 80'h0010ffabffabffabffab;
mem[7720] = 80'h0010ffabffabffabffab;
mem[7721] = 80'h0010ffabffabffabffab;
mem[7722] = 80'h0010ffabffabffabffab;
mem[7723] = 80'h0010ffabffabffabffab;
mem[7724] = 80'h0010ffabffabffabffab;
mem[7725] = 80'h0010ffabffabffabffab;
mem[7726] = 80'h0010ffabffabffabffab;
mem[7727] = 80'h0010ffabffabffabffab;
mem[7728] = 80'h0010ffabffabffabffab;
mem[7729] = 80'h0010ffabffabffabffab;
mem[7730] = 80'h0010ffabffabffabffab;
mem[7731] = 80'h0010ffabffabffabffab;
mem[7732] = 80'h0010ffabffabffabffab;
mem[7733] = 80'h0010ffabffabffabffab;
mem[7734] = 80'h0010ffabffabffabffab;
mem[7735] = 80'h0010ffabffabffabffab;
mem[7736] = 80'h0010ffabffabffabffab;
mem[7737] = 80'h0010ffabffabffabffab;
mem[7738] = 80'h0010ffabffabffabffab;
mem[7739] = 80'h0010ffabffabffabffab;
mem[7740] = 80'h0010ffabffabffabffab;
mem[7741] = 80'h0010ffabffabffabffab;
mem[7742] = 80'h0010ffabffabffabffab;
mem[7743] = 80'h0010ffabffabffabffab;
mem[7744] = 80'h0010ffabffabffabffab;
mem[7745] = 80'h0010ffabffabffabffab;
mem[7746] = 80'h0010ffabffabffabffab;
mem[7747] = 80'h0010ffabffabffabffab;
mem[7748] = 80'h0010ffabffabffabffab;
mem[7749] = 80'h0010ffabffabffabffab;
mem[7750] = 80'h0010ffabffabffabffab;
mem[7751] = 80'h0010ffabffabffabffab;
mem[7752] = 80'h0010ffabffabffabffab;
mem[7753] = 80'h0010ffabffabffabffab;
mem[7754] = 80'h0010ffabffabffabffab;
mem[7755] = 80'h0010ffabffabffabffab;
mem[7756] = 80'h0010ffabffabffabffab;
mem[7757] = 80'h0010ffabffabffabffab;
mem[7758] = 80'h0010ffabffabffabffab;
mem[7759] = 80'h0010ffabffabffabffab;
mem[7760] = 80'h0010ffabffabffabffab;
mem[7761] = 80'h0010ffabffabffabffab;
mem[7762] = 80'h0010ffabffabffabffab;
mem[7763] = 80'h0010ffabffabffabffab;
mem[7764] = 80'h0010ffabffabffabffab;
mem[7765] = 80'h0010ffabffabffabffab;
mem[7766] = 80'h0010ffabffabffabffab;
mem[7767] = 80'h0010ffabffabffabffab;
mem[7768] = 80'h0010ffabffabffabffab;
mem[7769] = 80'h0010ffabffabffabffab;
mem[7770] = 80'h0010ffabffabffabffab;
mem[7771] = 80'h0010ffabffabffabffab;
mem[7772] = 80'h0010ffabffabffabffab;
mem[7773] = 80'h0010ffabffabffabffab;
mem[7774] = 80'h0010ffabffabffabffab;
mem[7775] = 80'h0010ffabffabff171de3;
mem[7776] = 80'h0010cd8715a38acaa186;
mem[7777] = 80'h00101ab1608272cbfa89;
mem[7778] = 80'h0115ea5f9b5516000000;
mem[7779] = 80'h00000000000000000000;
mem[7780] = 80'h00000000000000000000;
mem[7781] = 80'h00000000000000000000;
mem[7782] = 80'h00000000000000000000;
mem[7783] = 80'h00000000000000000000;
mem[7784] = 80'h00000000000000000000;
mem[7785] = 80'h00000000000000000000;
mem[7786] = 80'h00000000000000000000;
mem[7787] = 80'h00000000000000000000;
mem[7788] = 80'h00000000000000000000;
mem[7789] = 80'h00000000000000000000;
mem[7790] = 80'h00000000000000000000;
mem[7791] = 80'h00000000000000000000;
mem[7792] = 80'h00000000000000000000;
mem[7793] = 80'h00000000000000000000;
mem[7794] = 80'h00000000000000000000;
mem[7795] = 80'h00000000000000000000;
mem[7796] = 80'h00000000000000000000;
mem[7797] = 80'h00000000000000000000;
mem[7798] = 80'h00000000000000000000;
mem[7799] = 80'h00000000000000000000;
mem[7800] = 80'h00000000000000000000;
mem[7801] = 80'h00000000000000000000;
mem[7802] = 80'h00000000000000000000;
mem[7803] = 80'h00000000000000000000;
mem[7804] = 80'h10100000010000010010;
mem[7805] = 80'h00109400000208004500;
mem[7806] = 80'h0010049089e90000fffd;
mem[7807] = 80'h0010ab2ec0550102c000;
mem[7808] = 80'h00100001ffabffabffab;
mem[7809] = 80'h0010ffabffabffabffab;
mem[7810] = 80'h0010ffabffabffabffab;
mem[7811] = 80'h0010ffabffabffabffab;
mem[7812] = 80'h0010ffabffabffabffab;
mem[7813] = 80'h0010ffabffabffabffab;
mem[7814] = 80'h0010ffabffabffabffab;
mem[7815] = 80'h0010ffabffabffabffab;
mem[7816] = 80'h0010ffabffabffabffab;
mem[7817] = 80'h0010ffabffabffabffab;
mem[7818] = 80'h0010ffabffabffabffab;
mem[7819] = 80'h0010ffabffabffabffab;
mem[7820] = 80'h0010ffabffabffabffab;
mem[7821] = 80'h0010ffabffabffabffab;
mem[7822] = 80'h0010ffabffabffabffab;
mem[7823] = 80'h0010ffabffabffabffab;
mem[7824] = 80'h0010ffabffabffabffab;
mem[7825] = 80'h0010ffabffabffabffab;
mem[7826] = 80'h0010ffabffabffabffab;
mem[7827] = 80'h0010ffabffabffabffab;
mem[7828] = 80'h0010ffabffabffabffab;
mem[7829] = 80'h0010ffabffabffabffab;
mem[7830] = 80'h0010ffabffabffabffab;
mem[7831] = 80'h0010ffabffabffabffab;
mem[7832] = 80'h0010ffabffabffabffab;
mem[7833] = 80'h0010ffabffabffabffab;
mem[7834] = 80'h0010ffabffabffabffab;
mem[7835] = 80'h0010ffabffabffabffab;
mem[7836] = 80'h0010ffabffabffabffab;
mem[7837] = 80'h0010ffabffabffabffab;
mem[7838] = 80'h0010ffabffabffabffab;
mem[7839] = 80'h0010ffabffabffabffab;
mem[7840] = 80'h0010ffabffabffabffab;
mem[7841] = 80'h0010ffabffabffabffab;
mem[7842] = 80'h0010ffabffabffabffab;
mem[7843] = 80'h0010ffabffabffabffab;
mem[7844] = 80'h0010ffabffabffabffab;
mem[7845] = 80'h0010ffabffabffabffab;
mem[7846] = 80'h0010ffabffabffabffab;
mem[7847] = 80'h0010ffabffabffabffab;
mem[7848] = 80'h0010ffabffabffabffab;
mem[7849] = 80'h0010ffabffabffabffab;
mem[7850] = 80'h0010ffabffabffabffab;
mem[7851] = 80'h0010ffabffabffabffab;
mem[7852] = 80'h0010ffabffabffabffab;
mem[7853] = 80'h0010ffabffabffabffab;
mem[7854] = 80'h0010ffabffabffabffab;
mem[7855] = 80'h0010ffabffabffabffab;
mem[7856] = 80'h0010ffabffabffabffab;
mem[7857] = 80'h0010ffabffabffabffab;
mem[7858] = 80'h0010ffabffabffabffab;
mem[7859] = 80'h0010ffabffabffabffab;
mem[7860] = 80'h0010ffabffabffabffab;
mem[7861] = 80'h0010ffabffabffabffab;
mem[7862] = 80'h0010ffabffabffabffab;
mem[7863] = 80'h0010ffabffabffabffab;
mem[7864] = 80'h0010ffabffabffabffab;
mem[7865] = 80'h0010ffabffabffabffab;
mem[7866] = 80'h0010ffabffabffabffab;
mem[7867] = 80'h0010ffabffabffabffab;
mem[7868] = 80'h0010ffabffabffabffab;
mem[7869] = 80'h0010ffabffabffabffab;
mem[7870] = 80'h0010ffabffabffabffab;
mem[7871] = 80'h0010ffabffabffabffab;
mem[7872] = 80'h0010ffabffabffabffab;
mem[7873] = 80'h0010ffabffabffabffab;
mem[7874] = 80'h0010ffabffabffabffab;
mem[7875] = 80'h0010ffabffabffabffab;
mem[7876] = 80'h0010ffabffabffabffab;
mem[7877] = 80'h0010ffabffabffabffab;
mem[7878] = 80'h0010ffabffabffabffab;
mem[7879] = 80'h0010ffabffabffabffab;
mem[7880] = 80'h0010ffabffabffabffab;
mem[7881] = 80'h0010ffabffabffabffab;
mem[7882] = 80'h0010ffabffabffabffab;
mem[7883] = 80'h0010ffabffabffabffab;
mem[7884] = 80'h0010ffabffabffabffab;
mem[7885] = 80'h0010ffabffabffabffab;
mem[7886] = 80'h0010ffabffabffabffab;
mem[7887] = 80'h0010ffabffabffabffab;
mem[7888] = 80'h0010ffabffabffabffab;
mem[7889] = 80'h0010ffabffabffabffab;
mem[7890] = 80'h0010ffabffabffabffab;
mem[7891] = 80'h0010ffabffabffabffab;
mem[7892] = 80'h0010ffabffabffabffab;
mem[7893] = 80'h0010ffabffabffabffab;
mem[7894] = 80'h0010ffabffabffabffab;
mem[7895] = 80'h0010ffabffabffabffab;
mem[7896] = 80'h0010ffabffabffabffab;
mem[7897] = 80'h0010ffabffabffabffab;
mem[7898] = 80'h0010ffabffabffabffab;
mem[7899] = 80'h0010ffabffabffabffab;
mem[7900] = 80'h0010ffabffabffabffab;
mem[7901] = 80'h0010ffabffabffabffab;
mem[7902] = 80'h0010ffabffabffabffab;
mem[7903] = 80'h0010ffabffabffabffab;
mem[7904] = 80'h0010ffabffabffabffab;
mem[7905] = 80'h0010ffabffabffabffab;
mem[7906] = 80'h0010ffabffabffabffab;
mem[7907] = 80'h0010ffabffabffabffab;
mem[7908] = 80'h0010ffabffabffabffab;
mem[7909] = 80'h0010ffabffabffabffab;
mem[7910] = 80'h0010ffabffabffabffab;
mem[7911] = 80'h0010ffabffabffabffab;
mem[7912] = 80'h0010ffabffabffabffab;
mem[7913] = 80'h0010ffabffabffabffab;
mem[7914] = 80'h0010ffabffabffabffab;
mem[7915] = 80'h0010ffabffabffabffab;
mem[7916] = 80'h0010ffabffabffabffab;
mem[7917] = 80'h0010ffabffabffabffab;
mem[7918] = 80'h0010ffabffabffabffab;
mem[7919] = 80'h0010ffabffabffabffab;
mem[7920] = 80'h0010ffabffabffabffab;
mem[7921] = 80'h0010ffabffabffabffab;
mem[7922] = 80'h0010ffabffabffabffab;
mem[7923] = 80'h0010ffabffabffabffab;
mem[7924] = 80'h0010ffabffabffabffab;
mem[7925] = 80'h0010ffabffabffabffab;
mem[7926] = 80'h0010ffabffabffabffab;
mem[7927] = 80'h0010ffabffabffabffab;
mem[7928] = 80'h0010ffabffabffabffab;
mem[7929] = 80'h0010ffabffabffabffab;
mem[7930] = 80'h0010ffabffabffabffab;
mem[7931] = 80'h0010ffabffabffabffab;
mem[7932] = 80'h0010ffabffabffabffab;
mem[7933] = 80'h0010ffabffabffabffab;
mem[7934] = 80'h0010ffabffabffabffab;
mem[7935] = 80'h0010ffabffabffabffab;
mem[7936] = 80'h0010ffabffabffabffab;
mem[7937] = 80'h0010ffabffabffabffab;
mem[7938] = 80'h0010ffabffabffabffab;
mem[7939] = 80'h0010ffabffabffabffab;
mem[7940] = 80'h0010ffabffabffabffab;
mem[7941] = 80'h0010ffabffabffabffab;
mem[7942] = 80'h0010ffabffabffabffab;
mem[7943] = 80'h0010ffabffabffabffab;
mem[7944] = 80'h0010ffabffabffabffab;
mem[7945] = 80'h0010ffabffabffabffab;
mem[7946] = 80'h0010ffabffabffabffab;
mem[7947] = 80'h0010ffabffabffabffab;
mem[7948] = 80'h0010ffabffabffabffab;
mem[7949] = 80'h0010ffab166c3de15f6c;
mem[7950] = 80'h00106135017301f744b1;
mem[7951] = 80'h0010c023e6aefc224668;
mem[7952] = 80'h011247b9000000000000;
mem[7953] = 80'h10100000010000010010;
mem[7954] = 80'h00109400000208004500;
mem[7955] = 80'h0010025f89ea0000fffd;
mem[7956] = 80'h0010ad5ec0550102c000;
mem[7957] = 80'h00100001ffabffabffab;
mem[7958] = 80'h0010ffabffabffabffab;
mem[7959] = 80'h0010ffabffabffabffab;
mem[7960] = 80'h0010ffabffabffabffab;
mem[7961] = 80'h0010ffabffabffabffab;
mem[7962] = 80'h0010ffabffabffabffab;
mem[7963] = 80'h0010ffabffabffabffab;
mem[7964] = 80'h0010ffabffabffabffab;
mem[7965] = 80'h0010ffabffabffabffab;
mem[7966] = 80'h0010ffabffabffabffab;
mem[7967] = 80'h0010ffabffabffabffab;
mem[7968] = 80'h0010ffabffabffabffab;
mem[7969] = 80'h0010ffabffabffabffab;
mem[7970] = 80'h0010ffabffabffabffab;
mem[7971] = 80'h0010ffabffabffabffab;
mem[7972] = 80'h0010ffabffabffabffab;
mem[7973] = 80'h0010ffabffabffabffab;
mem[7974] = 80'h0010ffabffabffabffab;
mem[7975] = 80'h0010ffabffabffabffab;
mem[7976] = 80'h0010ffabffabffabffab;
mem[7977] = 80'h0010ffabffabffabffab;
mem[7978] = 80'h0010ffabffabffabffab;
mem[7979] = 80'h0010ffabffabffabffab;
mem[7980] = 80'h0010ffabffabffabffab;
mem[7981] = 80'h0010ffabffabffabffab;
mem[7982] = 80'h0010ffabffabffabffab;
mem[7983] = 80'h0010ffabffabffabffab;
mem[7984] = 80'h0010ffabffabffabffab;
mem[7985] = 80'h0010ffabffabffabffab;
mem[7986] = 80'h0010ffabffabffabffab;
mem[7987] = 80'h0010ffabffabffabffab;
mem[7988] = 80'h0010ffabffabffabffab;
mem[7989] = 80'h0010ffabffabffabffab;
mem[7990] = 80'h0010ffabffabffabffab;
mem[7991] = 80'h0010ffabffabffabffab;
mem[7992] = 80'h0010ffabffabffabffab;
mem[7993] = 80'h0010ffabffabffabffab;
mem[7994] = 80'h0010ffabffabffabffab;
mem[7995] = 80'h0010ffabffabffabffab;
mem[7996] = 80'h0010ffabffabffabffab;
mem[7997] = 80'h0010ffabffabffabffab;
mem[7998] = 80'h0010ffabffabffabffab;
mem[7999] = 80'h0010ffabffabffabffab;
mem[8000] = 80'h0010ffabffabffabffab;
mem[8001] = 80'h0010ffabffabffabffab;
mem[8002] = 80'h0010ffabffabffabffab;
mem[8003] = 80'h0010ffabffabffabffab;
mem[8004] = 80'h0010ffabffabffabffab;
mem[8005] = 80'h0010ffabffabffabffab;
mem[8006] = 80'h0010ffabffabffabffab;
mem[8007] = 80'h0010ffabffabffabffab;
mem[8008] = 80'h0010ffabffabffabffab;
mem[8009] = 80'h0010ffabffabffabffab;
mem[8010] = 80'h0010ffabffabffabffab;
mem[8011] = 80'h0010ffabffabffabffab;
mem[8012] = 80'h0010ffabffabffabffab;
mem[8013] = 80'h0010ffabffabffabffab;
mem[8014] = 80'h0010ffabffabffabffab;
mem[8015] = 80'h0010ffabffabffabffab;
mem[8016] = 80'h0010ffabffabffabffab;
mem[8017] = 80'h0010ffabffabffabffab;
mem[8018] = 80'h0010ffabffabffabffab;
mem[8019] = 80'h0010ffabffabffabffab;
mem[8020] = 80'h0010ffabffabffabffab;
mem[8021] = 80'h0010ffabffabffabffab;
mem[8022] = 80'h0010ffabffabffabffab;
mem[8023] = 80'h0010ffabffabffabffab;
mem[8024] = 80'h0010ffabffabffabffab;
mem[8025] = 80'h0010ffabffabffabffab;
mem[8026] = 80'h0010ffabffabffabffab;
mem[8027] = 80'h0010ffabffabffabffab;
mem[8028] = 80'h0010ff15fe5f9437e626;
mem[8029] = 80'h0010f55d0489c15acfed;
mem[8030] = 80'h0010d10f6aecc09f874a;
mem[8031] = 80'h01118c00000000000000;
mem[8032] = 80'h10100000010000010010;
mem[8033] = 80'h00109400000208004500;
mem[8034] = 80'h0010014589eb0000fffd;
mem[8035] = 80'h0010ae77c0550102c000;
mem[8036] = 80'h00100001ffabffabffab;
mem[8037] = 80'h0010ffabffabffabffab;
mem[8038] = 80'h0010ffabffabffabffab;
mem[8039] = 80'h0010ffabffabffabffab;
mem[8040] = 80'h0010ffabffabffabffab;
mem[8041] = 80'h0010ffabffabffabffab;
mem[8042] = 80'h0010ffabffabffabffab;
mem[8043] = 80'h0010ffabffabffabffab;
mem[8044] = 80'h0010ffabffabffabffab;
mem[8045] = 80'h0010ffabffabffabffab;
mem[8046] = 80'h0010ffabffabffabffab;
mem[8047] = 80'h0010ffabffabffabffab;
mem[8048] = 80'h0010ffabffabffabffab;
mem[8049] = 80'h0010ffabffabffabffab;
mem[8050] = 80'h0010ffabffabffabffab;
mem[8051] = 80'h0010ffabffabffabffab;
mem[8052] = 80'h0010ffabffabffabffab;
mem[8053] = 80'h0010ffabffabffabffab;
mem[8054] = 80'h0010ffabffabffabffab;
mem[8055] = 80'h0010ffabffabffabffab;
mem[8056] = 80'h0010ffabffabffabffab;
mem[8057] = 80'h0010ffabffabffabffab;
mem[8058] = 80'h0010ffabffabffabffab;
mem[8059] = 80'h0010ffabffabffabffab;
mem[8060] = 80'h0010ffabffabffabffab;
mem[8061] = 80'h0010ffabffabffabffab;
mem[8062] = 80'h0010ffabffabffabffab;
mem[8063] = 80'h0010ffabffabffabffab;
mem[8064] = 80'h0010ffabffabffabffab;
mem[8065] = 80'h0010ffabffabffabffab;
mem[8066] = 80'h0010ffabffabffabffab;
mem[8067] = 80'h0010ffabffabffabffab;
mem[8068] = 80'h0010ffabffabffabffab;
mem[8069] = 80'h0010ffabffabffabffab;
mem[8070] = 80'h0010ffabffabffabffab;
mem[8071] = 80'h0010ffabffabffabff14;
mem[8072] = 80'h00108f81b8ef9fe44a96;
mem[8073] = 80'h0010d60e2caf1cb880d6;
mem[8074] = 80'h0117bab272f5f10b2a00;
mem[8075] = 80'h00000000000000000000;
mem[8076] = 80'h00000000000000000000;
mem[8077] = 80'h00000000000000000000;
mem[8078] = 80'h00000000000000000000;
mem[8079] = 80'h00000000000000000000;
mem[8080] = 80'h00000000000000000000;
mem[8081] = 80'h00000000000000000000;
mem[8082] = 80'h00000000000000000000;
mem[8083] = 80'h00000000000000000000;
mem[8084] = 80'h00000000000000000000;
mem[8085] = 80'h00000000000000000000;
mem[8086] = 80'h00000000000000000000;
mem[8087] = 80'h00000000000000000000;
mem[8088] = 80'h00000000000000000000;
mem[8089] = 80'h00000000000000000000;
mem[8090] = 80'h00000000000000000000;
mem[8091] = 80'h00000000000000000000;
mem[8092] = 80'h00000000000000000000;
mem[8093] = 80'h00000000000000000000;
mem[8094] = 80'h00000000000000000000;
mem[8095] = 80'h00000000000000000000;
mem[8096] = 80'h00000000000000000000;
mem[8097] = 80'h00000000000000000000;
mem[8098] = 80'h00000000000000000000;
mem[8099] = 80'h00000000000000000000;
mem[8100] = 80'h00000000000000000000;
mem[8101] = 80'h00000000000000000000;
mem[8102] = 80'h00000000000000000000;
mem[8103] = 80'h00000000000000000000;
mem[8104] = 80'h00000000000000000000;
mem[8105] = 80'h00000000000000000000;
mem[8106] = 80'h00000000000000000000;
mem[8107] = 80'h00000000000000000000;
mem[8108] = 80'h00000000000000000000;
mem[8109] = 80'h00000000000000000000;
mem[8110] = 80'h00000000000000000000;
mem[8111] = 80'h00000000000000000000;
mem[8112] = 80'h00000000000000000000;
mem[8113] = 80'h00000000000000000000;
mem[8114] = 80'h00000000000000000000;
mem[8115] = 80'h00000000000000000000;
mem[8116] = 80'h00000000000000000000;
mem[8117] = 80'h00000000000000000000;
mem[8118] = 80'h00000000000000000000;
mem[8119] = 80'h00000000000000000000;
mem[8120] = 80'h00000000000000000000;
mem[8121] = 80'h00000000000000000000;
mem[8122] = 80'h00000000000000000000;
mem[8123] = 80'h00000000000000000000;
mem[8124] = 80'h00000000000000000000;
mem[8125] = 80'h00000000000000000000;
mem[8126] = 80'h00000000000000000000;
mem[8127] = 80'h00000000000000000000;
mem[8128] = 80'h00000000000000000000;
mem[8129] = 80'h00000000000000000000;
mem[8130] = 80'h00000000000000000000;
mem[8131] = 80'h00000000000000000000;
mem[8132] = 80'h00000000000000000000;
mem[8133] = 80'h00000000000000000000;
mem[8134] = 80'h00000000000000000000;
mem[8135] = 80'h00000000000000000000;
mem[8136] = 80'h00000000000000000000;
mem[8137] = 80'h00000000000000000000;
mem[8138] = 80'h00000000000000000000;
mem[8139] = 80'h00000000000000000000;
mem[8140] = 80'h00000000000000000000;
mem[8141] = 80'h00000000000000000000;
mem[8142] = 80'h00000000000000000000;
mem[8143] = 80'h00000000000000000000;
mem[8144] = 80'h00000000000000000000;
mem[8145] = 80'h00000000000000000000;
mem[8146] = 80'h00000000000000000000;
mem[8147] = 80'h00000000000000000000;
mem[8148] = 80'h00000000000000000000;
mem[8149] = 80'h00000000000000000000;
mem[8150] = 80'h00000000000000000000;
mem[8151] = 80'h00000000000000000000;
mem[8152] = 80'h00000000000000000000;
mem[8153] = 80'h00000000000000000000;
mem[8154] = 80'h00000000000000000000;
mem[8155] = 80'h00000000000000000000;
mem[8156] = 80'h00000000000000000000;
mem[8157] = 80'h00000000000000000000;
mem[8158] = 80'h00000000000000000000;
mem[8159] = 80'h00000000000000000000;
mem[8160] = 80'h00000000000000000000;
mem[8161] = 80'h00000000000000000000;
mem[8162] = 80'h00000000000000000000;
mem[8163] = 80'h00000000000000000000;
mem[8164] = 80'h00000000000000000000;
mem[8165] = 80'h00000000000000000000;
mem[8166] = 80'h00000000000000000000;
mem[8167] = 80'h00000000000000000000;
mem[8168] = 80'h00000000000000000000;
mem[8169] = 80'h00000000000000000000;
mem[8170] = 80'h00000000000000000000;
mem[8171] = 80'h00000000000000000000;
mem[8172] = 80'h00000000000000000000;
mem[8173] = 80'h00000000000000000000;
mem[8174] = 80'h00000000000000000000;
mem[8175] = 80'h00000000000000000000;
mem[8176] = 80'h00000000000000000000;
mem[8177] = 80'h00000000000000000000;
mem[8178] = 80'h00000000000000000000;
mem[8179] = 80'h00000000000000000000;
mem[8180] = 80'h00000000000000000000;
mem[8181] = 80'h00000000000000000000;
mem[8182] = 80'h00000000000000000000;
mem[8183] = 80'h00000000000000000000;
mem[8184] = 80'h00000000000000000000;
mem[8185] = 80'h00000000000000000000;
mem[8186] = 80'h00000000000000000000;
mem[8187] = 80'h00000000000000000000;
mem[8188] = 80'h00000000000000000000;
mem[8189] = 80'h00000000000000000000;
mem[8190] = 80'h00000000000000000000;
mem[8191] = 80'h00000000000000000000;
end


//*********************
//MAIN CORE
//********************* 
reg [15:0] time_cnt ;    
reg [31:0] cnt ;

initial begin
    time_cnt = 'd0 ;
    cnt      = 'd0 ;
end

always @(posedge clk) begin

    if ( time_cnt == 'd1000 ) begin
        time_cnt <= time_cnt ;
    end
    else begin
        time_cnt <= time_cnt+1'b1 ;
    end
end

always @(posedge clk) begin

    if ( time_cnt >'d900 ) begin
        if ( cnt == 'd8191 ) begin
            cnt <= 'd0 ;
        end
        else begin
           cnt <= cnt+1'b1 ; 
        end
    end
    else begin
        cnt <= 'd0 ;
    end
end

wire [12:0] rd_addr ;

assign rd_addr = cnt[12:0] ;


always @(posedge clk) begin
	dout_ff <= mem[rd_addr] ;
end


assign sop  = dout_ff[76] ;
assign eop  = dout_ff[72] ;
assign dval = dout_ff[68] ;
assign mod  = dout_ff[66:64] ;
assign dout = dout_ff[63:0] ;


//*********************
endmodule   