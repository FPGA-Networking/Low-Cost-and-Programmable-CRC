

// **************************************************************
// COPYRIGHT(c)2015, Xidian University
// All rights reserved.
//
// IP LIB INDEX :  
// IP Name      :      
// File name    : 
// Module name  : 
// Full name    :  
//
// Author       : Liu-Huan 
// Email        : assasin9997@163.com 
// Data         : 
// Version      : V 1.0 
// 
// Abstract     : 
// Called by    :  
// 
// Modification history
// -----------------------------------------------------------------
// 
// 
//
// *****************************************************************

// *******************
// TIMESCALE
// ******************* 
`timescale 1ns/1ps 

// *******************
// INFORMATION
// *******************


//*******************
//DEFINE(s)
//*******************
//`define UDLY 1    //Unit delay, for non-blocking assignments in sequential logic



//*******************
//DEFINE MODULE PORT
//*******************
module  go_ahead_4096

# ( parameter  [1023:0] AHEAD_POLY = 0 )


 (     
        input           clk ,
        input           rst ,

        input           crc_en_i,
        input   [31:0]  crc_i,  
        output reg         crc_en_o,
        output reg [31:0]  crc_o


              ) ;

//*******************
//DEFINE LOCAL PARAMETER
//*******************
//parameter(s)
 





// reg [1023:0] ahead = AHEAD_POLY ;
// wire [8:0] test ;

wire [31:0] ahead ;






















//*********************
//INNER SIGNAL DECLARATION
//*********************

 
// crc-32
  //   function [31:0] CRC32_ahead;

  //   input [31:0] crc_i;
  //   // input [31:0] crc_o;
  //   //reg [31:0] d;
  //   reg [31:0] c;
  //   reg [31:0] newcrc;
  // begin
  //   c = crc_i;

  //   newcrc[0 ]  = (c[0]&AHEAD_POLY[1023-32* 0  ])^(c[1]&AHEAD_POLY[1023-32* 0  -1])^(c[2]&AHEAD_POLY[1023-32* -2 ])^(c[3]&AHEAD_POLY[1023-32* 0  -3])^(c[4]&AHEAD_POLY[1023-32* 0  -4])^(c[5]&AHEAD_POLY[1023-32* 0  -5])^(c[6]&AHEAD_POLY[1023-32* 0  -6])^(c[7]&AHEAD_POLY[1023-32* 0  -7])^(c[8]&AHEAD_POLY[1023-32* 0  -8])^(c[9]&AHEAD_POLY[1023-32* 0  -9])^(c[10]&AHEAD_POLY[1023-32* 0  -10])^(c[11]&AHEAD_POLY[1023-32* 0  -11])^(c[12]&AHEAD_POLY[1023-32* 0  -12])^(c[13]&AHEAD_POLY[1023-32* 0  -13])^(c[14]&AHEAD_POLY[1023-32* 0  -14])^(c[15]&AHEAD_POLY[1023-32* 0  -15])^(c[16]&AHEAD_POLY[1023-32* 0  -16])^(c[17]&AHEAD_POLY[1023-32* 0  -17])^(c[18]&AHEAD_POLY[1023-32* 0  -18])^(c[19]&AHEAD_POLY[1023-32* 0  -19])^(c[20]&AHEAD_POLY[1023-32* 0  -20])^(c[21]&AHEAD_POLY[1023-32* 0  -21])^(c[22]&AHEAD_POLY[1023-32* 0  -22])^(c[23]&AHEAD_POLY[1023-32* 0  -23])^(c[24]&AHEAD_POLY[1023-32* 0  -24])^(c[25]&AHEAD_POLY[1023-32* 0  -25])^(c[26]&AHEAD_POLY[1023-32* 0  -26])^(c[27]&AHEAD_POLY[1023-32* 0  -27])^(c[28]&AHEAD_POLY[1023-32* 0  -28])^(c[29]&AHEAD_POLY[1023-32* 0  -29])^(c[30]&AHEAD_POLY[1023-32* 0  -30])^(c[31]&AHEAD_POLY[1023-32* 0  -31]);
  //   newcrc[1 ]  = (c[0]&AHEAD_POLY[1023-32* 1  ])^(c[1]&AHEAD_POLY[1023-32* 1  -1])^(c[2]&AHEAD_POLY[1023-32* -2 ])^(c[3]&AHEAD_POLY[1023-32* 1  -3])^(c[4]&AHEAD_POLY[1023-32* 1  -4])^(c[5]&AHEAD_POLY[1023-32* 1  -5])^(c[6]&AHEAD_POLY[1023-32* 1  -6])^(c[7]&AHEAD_POLY[1023-32* 1  -7])^(c[8]&AHEAD_POLY[1023-32* 1  -8])^(c[9]&AHEAD_POLY[1023-32* 1  -9])^(c[10]&AHEAD_POLY[1023-32* 1  -10])^(c[11]&AHEAD_POLY[1023-32* 1  -11])^(c[12]&AHEAD_POLY[1023-32* 1  -12])^(c[13]&AHEAD_POLY[1023-32* 1  -13])^(c[14]&AHEAD_POLY[1023-32* 1  -14])^(c[15]&AHEAD_POLY[1023-32* 1  -15])^(c[16]&AHEAD_POLY[1023-32* 1  -16])^(c[17]&AHEAD_POLY[1023-32* 1  -17])^(c[18]&AHEAD_POLY[1023-32* 1  -18])^(c[19]&AHEAD_POLY[1023-32* 1  -19])^(c[20]&AHEAD_POLY[1023-32* 1  -20])^(c[21]&AHEAD_POLY[1023-32* 1  -21])^(c[22]&AHEAD_POLY[1023-32* 1  -22])^(c[23]&AHEAD_POLY[1023-32* 1  -23])^(c[24]&AHEAD_POLY[1023-32* 1  -24])^(c[25]&AHEAD_POLY[1023-32* 1  -25])^(c[26]&AHEAD_POLY[1023-32* 1  -26])^(c[27]&AHEAD_POLY[1023-32* 1  -27])^(c[28]&AHEAD_POLY[1023-32* 1  -28])^(c[29]&AHEAD_POLY[1023-32* 1  -29])^(c[30]&AHEAD_POLY[1023-32* 1  -30])^(c[31]&AHEAD_POLY[1023-32* 1  -31]);
  //   newcrc[2 ]  = (c[0]&AHEAD_POLY[1023-32* 2  ])^(c[1]&AHEAD_POLY[1023-32* 2  -1])^(c[2]&AHEAD_POLY[1023-32* -2 ])^(c[3]&AHEAD_POLY[1023-32* 2  -3])^(c[4]&AHEAD_POLY[1023-32* 2  -4])^(c[5]&AHEAD_POLY[1023-32* 2  -5])^(c[6]&AHEAD_POLY[1023-32* 2  -6])^(c[7]&AHEAD_POLY[1023-32* 2  -7])^(c[8]&AHEAD_POLY[1023-32* 2  -8])^(c[9]&AHEAD_POLY[1023-32* 2  -9])^(c[10]&AHEAD_POLY[1023-32* 2  -10])^(c[11]&AHEAD_POLY[1023-32* 2  -11])^(c[12]&AHEAD_POLY[1023-32* 2  -12])^(c[13]&AHEAD_POLY[1023-32* 2  -13])^(c[14]&AHEAD_POLY[1023-32* 2  -14])^(c[15]&AHEAD_POLY[1023-32* 2  -15])^(c[16]&AHEAD_POLY[1023-32* 2  -16])^(c[17]&AHEAD_POLY[1023-32* 2  -17])^(c[18]&AHEAD_POLY[1023-32* 2  -18])^(c[19]&AHEAD_POLY[1023-32* 2  -19])^(c[20]&AHEAD_POLY[1023-32* 2  -20])^(c[21]&AHEAD_POLY[1023-32* 2  -21])^(c[22]&AHEAD_POLY[1023-32* 2  -22])^(c[23]&AHEAD_POLY[1023-32* 2  -23])^(c[24]&AHEAD_POLY[1023-32* 2  -24])^(c[25]&AHEAD_POLY[1023-32* 2  -25])^(c[26]&AHEAD_POLY[1023-32* 2  -26])^(c[27]&AHEAD_POLY[1023-32* 2  -27])^(c[28]&AHEAD_POLY[1023-32* 2  -28])^(c[29]&AHEAD_POLY[1023-32* 2  -29])^(c[30]&AHEAD_POLY[1023-32* 2  -30])^(c[31]&AHEAD_POLY[1023-32* 2  -31]);
  //   newcrc[3 ]  = (c[0]&AHEAD_POLY[1023-32* 3  ])^(c[1]&AHEAD_POLY[1023-32* 3  -1])^(c[2]&AHEAD_POLY[1023-32* -2 ])^(c[3]&AHEAD_POLY[1023-32* 3  -3])^(c[4]&AHEAD_POLY[1023-32* 3  -4])^(c[5]&AHEAD_POLY[1023-32* 3  -5])^(c[6]&AHEAD_POLY[1023-32* 3  -6])^(c[7]&AHEAD_POLY[1023-32* 3  -7])^(c[8]&AHEAD_POLY[1023-32* 3  -8])^(c[9]&AHEAD_POLY[1023-32* 3  -9])^(c[10]&AHEAD_POLY[1023-32* 3  -10])^(c[11]&AHEAD_POLY[1023-32* 3  -11])^(c[12]&AHEAD_POLY[1023-32* 3  -12])^(c[13]&AHEAD_POLY[1023-32* 3  -13])^(c[14]&AHEAD_POLY[1023-32* 3  -14])^(c[15]&AHEAD_POLY[1023-32* 3  -15])^(c[16]&AHEAD_POLY[1023-32* 3  -16])^(c[17]&AHEAD_POLY[1023-32* 3  -17])^(c[18]&AHEAD_POLY[1023-32* 3  -18])^(c[19]&AHEAD_POLY[1023-32* 3  -19])^(c[20]&AHEAD_POLY[1023-32* 3  -20])^(c[21]&AHEAD_POLY[1023-32* 3  -21])^(c[22]&AHEAD_POLY[1023-32* 3  -22])^(c[23]&AHEAD_POLY[1023-32* 3  -23])^(c[24]&AHEAD_POLY[1023-32* 3  -24])^(c[25]&AHEAD_POLY[1023-32* 3  -25])^(c[26]&AHEAD_POLY[1023-32* 3  -26])^(c[27]&AHEAD_POLY[1023-32* 3  -27])^(c[28]&AHEAD_POLY[1023-32* 3  -28])^(c[29]&AHEAD_POLY[1023-32* 3  -29])^(c[30]&AHEAD_POLY[1023-32* 3  -30])^(c[31]&AHEAD_POLY[1023-32* 3  -31]);
  //   newcrc[4 ]  = (c[0]&AHEAD_POLY[1023-32* 4  ])^(c[1]&AHEAD_POLY[1023-32* 4  -1])^(c[2]&AHEAD_POLY[1023-32* -2 ])^(c[3]&AHEAD_POLY[1023-32* 4  -3])^(c[4]&AHEAD_POLY[1023-32* 4  -4])^(c[5]&AHEAD_POLY[1023-32* 4  -5])^(c[6]&AHEAD_POLY[1023-32* 4  -6])^(c[7]&AHEAD_POLY[1023-32* 4  -7])^(c[8]&AHEAD_POLY[1023-32* 4  -8])^(c[9]&AHEAD_POLY[1023-32* 4  -9])^(c[10]&AHEAD_POLY[1023-32* 4  -10])^(c[11]&AHEAD_POLY[1023-32* 4  -11])^(c[12]&AHEAD_POLY[1023-32* 4  -12])^(c[13]&AHEAD_POLY[1023-32* 4  -13])^(c[14]&AHEAD_POLY[1023-32* 4  -14])^(c[15]&AHEAD_POLY[1023-32* 4  -15])^(c[16]&AHEAD_POLY[1023-32* 4  -16])^(c[17]&AHEAD_POLY[1023-32* 4  -17])^(c[18]&AHEAD_POLY[1023-32* 4  -18])^(c[19]&AHEAD_POLY[1023-32* 4  -19])^(c[20]&AHEAD_POLY[1023-32* 4  -20])^(c[21]&AHEAD_POLY[1023-32* 4  -21])^(c[22]&AHEAD_POLY[1023-32* 4  -22])^(c[23]&AHEAD_POLY[1023-32* 4  -23])^(c[24]&AHEAD_POLY[1023-32* 4  -24])^(c[25]&AHEAD_POLY[1023-32* 4  -25])^(c[26]&AHEAD_POLY[1023-32* 4  -26])^(c[27]&AHEAD_POLY[1023-32* 4  -27])^(c[28]&AHEAD_POLY[1023-32* 4  -28])^(c[29]&AHEAD_POLY[1023-32* 4  -29])^(c[30]&AHEAD_POLY[1023-32* 4  -30])^(c[31]&AHEAD_POLY[1023-32* 4  -31]);
  //   newcrc[5 ]  = (c[0]&AHEAD_POLY[1023-32* 5  ])^(c[1]&AHEAD_POLY[1023-32* 5  -1])^(c[2]&AHEAD_POLY[1023-32* -2 ])^(c[3]&AHEAD_POLY[1023-32* 5  -3])^(c[4]&AHEAD_POLY[1023-32* 5  -4])^(c[5]&AHEAD_POLY[1023-32* 5  -5])^(c[6]&AHEAD_POLY[1023-32* 5  -6])^(c[7]&AHEAD_POLY[1023-32* 5  -7])^(c[8]&AHEAD_POLY[1023-32* 5  -8])^(c[9]&AHEAD_POLY[1023-32* 5  -9])^(c[10]&AHEAD_POLY[1023-32* 5  -10])^(c[11]&AHEAD_POLY[1023-32* 5  -11])^(c[12]&AHEAD_POLY[1023-32* 5  -12])^(c[13]&AHEAD_POLY[1023-32* 5  -13])^(c[14]&AHEAD_POLY[1023-32* 5  -14])^(c[15]&AHEAD_POLY[1023-32* 5  -15])^(c[16]&AHEAD_POLY[1023-32* 5  -16])^(c[17]&AHEAD_POLY[1023-32* 5  -17])^(c[18]&AHEAD_POLY[1023-32* 5  -18])^(c[19]&AHEAD_POLY[1023-32* 5  -19])^(c[20]&AHEAD_POLY[1023-32* 5  -20])^(c[21]&AHEAD_POLY[1023-32* 5  -21])^(c[22]&AHEAD_POLY[1023-32* 5  -22])^(c[23]&AHEAD_POLY[1023-32* 5  -23])^(c[24]&AHEAD_POLY[1023-32* 5  -24])^(c[25]&AHEAD_POLY[1023-32* 5  -25])^(c[26]&AHEAD_POLY[1023-32* 5  -26])^(c[27]&AHEAD_POLY[1023-32* 5  -27])^(c[28]&AHEAD_POLY[1023-32* 5  -28])^(c[29]&AHEAD_POLY[1023-32* 5  -29])^(c[30]&AHEAD_POLY[1023-32* 5  -30])^(c[31]&AHEAD_POLY[1023-32* 5  -31]);
  //   newcrc[6 ]  = (c[0]&AHEAD_POLY[1023-32* 6  ])^(c[1]&AHEAD_POLY[1023-32* 6  -1])^(c[2]&AHEAD_POLY[1023-32* -2 ])^(c[3]&AHEAD_POLY[1023-32* 6  -3])^(c[4]&AHEAD_POLY[1023-32* 6  -4])^(c[5]&AHEAD_POLY[1023-32* 6  -5])^(c[6]&AHEAD_POLY[1023-32* 6  -6])^(c[7]&AHEAD_POLY[1023-32* 6  -7])^(c[8]&AHEAD_POLY[1023-32* 6  -8])^(c[9]&AHEAD_POLY[1023-32* 6  -9])^(c[10]&AHEAD_POLY[1023-32* 6  -10])^(c[11]&AHEAD_POLY[1023-32* 6  -11])^(c[12]&AHEAD_POLY[1023-32* 6  -12])^(c[13]&AHEAD_POLY[1023-32* 6  -13])^(c[14]&AHEAD_POLY[1023-32* 6  -14])^(c[15]&AHEAD_POLY[1023-32* 6  -15])^(c[16]&AHEAD_POLY[1023-32* 6  -16])^(c[17]&AHEAD_POLY[1023-32* 6  -17])^(c[18]&AHEAD_POLY[1023-32* 6  -18])^(c[19]&AHEAD_POLY[1023-32* 6  -19])^(c[20]&AHEAD_POLY[1023-32* 6  -20])^(c[21]&AHEAD_POLY[1023-32* 6  -21])^(c[22]&AHEAD_POLY[1023-32* 6  -22])^(c[23]&AHEAD_POLY[1023-32* 6  -23])^(c[24]&AHEAD_POLY[1023-32* 6  -24])^(c[25]&AHEAD_POLY[1023-32* 6  -25])^(c[26]&AHEAD_POLY[1023-32* 6  -26])^(c[27]&AHEAD_POLY[1023-32* 6  -27])^(c[28]&AHEAD_POLY[1023-32* 6  -28])^(c[29]&AHEAD_POLY[1023-32* 6  -29])^(c[30]&AHEAD_POLY[1023-32* 6  -30])^(c[31]&AHEAD_POLY[1023-32* 6  -31]);
  //   newcrc[7 ]  = (c[0]&AHEAD_POLY[1023-32* 7  ])^(c[1]&AHEAD_POLY[1023-32* 7  -1])^(c[2]&AHEAD_POLY[1023-32* -2 ])^(c[3]&AHEAD_POLY[1023-32* 7  -3])^(c[4]&AHEAD_POLY[1023-32* 7  -4])^(c[5]&AHEAD_POLY[1023-32* 7  -5])^(c[6]&AHEAD_POLY[1023-32* 7  -6])^(c[7]&AHEAD_POLY[1023-32* 7  -7])^(c[8]&AHEAD_POLY[1023-32* 7  -8])^(c[9]&AHEAD_POLY[1023-32* 7  -9])^(c[10]&AHEAD_POLY[1023-32* 7  -10])^(c[11]&AHEAD_POLY[1023-32* 7  -11])^(c[12]&AHEAD_POLY[1023-32* 7  -12])^(c[13]&AHEAD_POLY[1023-32* 7  -13])^(c[14]&AHEAD_POLY[1023-32* 7  -14])^(c[15]&AHEAD_POLY[1023-32* 7  -15])^(c[16]&AHEAD_POLY[1023-32* 7  -16])^(c[17]&AHEAD_POLY[1023-32* 7  -17])^(c[18]&AHEAD_POLY[1023-32* 7  -18])^(c[19]&AHEAD_POLY[1023-32* 7  -19])^(c[20]&AHEAD_POLY[1023-32* 7  -20])^(c[21]&AHEAD_POLY[1023-32* 7  -21])^(c[22]&AHEAD_POLY[1023-32* 7  -22])^(c[23]&AHEAD_POLY[1023-32* 7  -23])^(c[24]&AHEAD_POLY[1023-32* 7  -24])^(c[25]&AHEAD_POLY[1023-32* 7  -25])^(c[26]&AHEAD_POLY[1023-32* 7  -26])^(c[27]&AHEAD_POLY[1023-32* 7  -27])^(c[28]&AHEAD_POLY[1023-32* 7  -28])^(c[29]&AHEAD_POLY[1023-32* 7  -29])^(c[30]&AHEAD_POLY[1023-32* 7  -30])^(c[31]&AHEAD_POLY[1023-32* 7  -31]);
  //   newcrc[8 ]  = (c[0]&AHEAD_POLY[1023-32* 8  ])^(c[1]&AHEAD_POLY[1023-32* 8  -1])^(c[2]&AHEAD_POLY[1023-32* -2 ])^(c[3]&AHEAD_POLY[1023-32* 8  -3])^(c[4]&AHEAD_POLY[1023-32* 8  -4])^(c[5]&AHEAD_POLY[1023-32* 8  -5])^(c[6]&AHEAD_POLY[1023-32* 8  -6])^(c[7]&AHEAD_POLY[1023-32* 8  -7])^(c[8]&AHEAD_POLY[1023-32* 8  -8])^(c[9]&AHEAD_POLY[1023-32* 8  -9])^(c[10]&AHEAD_POLY[1023-32* 8  -10])^(c[11]&AHEAD_POLY[1023-32* 8  -11])^(c[12]&AHEAD_POLY[1023-32* 8  -12])^(c[13]&AHEAD_POLY[1023-32* 8  -13])^(c[14]&AHEAD_POLY[1023-32* 8  -14])^(c[15]&AHEAD_POLY[1023-32* 8  -15])^(c[16]&AHEAD_POLY[1023-32* 8  -16])^(c[17]&AHEAD_POLY[1023-32* 8  -17])^(c[18]&AHEAD_POLY[1023-32* 8  -18])^(c[19]&AHEAD_POLY[1023-32* 8  -19])^(c[20]&AHEAD_POLY[1023-32* 8  -20])^(c[21]&AHEAD_POLY[1023-32* 8  -21])^(c[22]&AHEAD_POLY[1023-32* 8  -22])^(c[23]&AHEAD_POLY[1023-32* 8  -23])^(c[24]&AHEAD_POLY[1023-32* 8  -24])^(c[25]&AHEAD_POLY[1023-32* 8  -25])^(c[26]&AHEAD_POLY[1023-32* 8  -26])^(c[27]&AHEAD_POLY[1023-32* 8  -27])^(c[28]&AHEAD_POLY[1023-32* 8  -28])^(c[29]&AHEAD_POLY[1023-32* 8  -29])^(c[30]&AHEAD_POLY[1023-32* 8  -30])^(c[31]&AHEAD_POLY[1023-32* 8  -31]);
  //   newcrc[9 ]  = (c[0]&AHEAD_POLY[1023-32* 9  ])^(c[1]&AHEAD_POLY[1023-32* 9  -1])^(c[2]&AHEAD_POLY[1023-32* -2 ])^(c[3]&AHEAD_POLY[1023-32* 9  -3])^(c[4]&AHEAD_POLY[1023-32* 9  -4])^(c[5]&AHEAD_POLY[1023-32* 9  -5])^(c[6]&AHEAD_POLY[1023-32* 9  -6])^(c[7]&AHEAD_POLY[1023-32* 9  -7])^(c[8]&AHEAD_POLY[1023-32* 9  -8])^(c[9]&AHEAD_POLY[1023-32* 9  -9])^(c[10]&AHEAD_POLY[1023-32* 9  -10])^(c[11]&AHEAD_POLY[1023-32* 9  -11])^(c[12]&AHEAD_POLY[1023-32* 9  -12])^(c[13]&AHEAD_POLY[1023-32* 9  -13])^(c[14]&AHEAD_POLY[1023-32* 9  -14])^(c[15]&AHEAD_POLY[1023-32* 9  -15])^(c[16]&AHEAD_POLY[1023-32* 9  -16])^(c[17]&AHEAD_POLY[1023-32* 9  -17])^(c[18]&AHEAD_POLY[1023-32* 9  -18])^(c[19]&AHEAD_POLY[1023-32* 9  -19])^(c[20]&AHEAD_POLY[1023-32* 9  -20])^(c[21]&AHEAD_POLY[1023-32* 9  -21])^(c[22]&AHEAD_POLY[1023-32* 9  -22])^(c[23]&AHEAD_POLY[1023-32* 9  -23])^(c[24]&AHEAD_POLY[1023-32* 9  -24])^(c[25]&AHEAD_POLY[1023-32* 9  -25])^(c[26]&AHEAD_POLY[1023-32* 9  -26])^(c[27]&AHEAD_POLY[1023-32* 9  -27])^(c[28]&AHEAD_POLY[1023-32* 9  -28])^(c[29]&AHEAD_POLY[1023-32* 9  -29])^(c[30]&AHEAD_POLY[1023-32* 9  -30])^(c[31]&AHEAD_POLY[1023-32* 9  -31]);
  //   newcrc[10]  = (c[0]&AHEAD_POLY[1023-32* 10 ])^(c[1]&AHEAD_POLY[1023-32* 10 -1])^(c[2]&AHEAD_POLY[1023-32* -2 ])^(c[3]&AHEAD_POLY[1023-32* 10 -3])^(c[4]&AHEAD_POLY[1023-32* 10 -4])^(c[5]&AHEAD_POLY[1023-32* 10 -5])^(c[6]&AHEAD_POLY[1023-32* 10 -6])^(c[7]&AHEAD_POLY[1023-32* 10 -7])^(c[8]&AHEAD_POLY[1023-32* 10 -8])^(c[9]&AHEAD_POLY[1023-32* 10 -9])^(c[10]&AHEAD_POLY[1023-32* 10 -10])^(c[11]&AHEAD_POLY[1023-32* 10 -11])^(c[12]&AHEAD_POLY[1023-32* 10 -12])^(c[13]&AHEAD_POLY[1023-32* 10 -13])^(c[14]&AHEAD_POLY[1023-32* 10 -14])^(c[15]&AHEAD_POLY[1023-32* 10 -15])^(c[16]&AHEAD_POLY[1023-32* 10 -16])^(c[17]&AHEAD_POLY[1023-32* 10 -17])^(c[18]&AHEAD_POLY[1023-32* 10 -18])^(c[19]&AHEAD_POLY[1023-32* 10 -19])^(c[20]&AHEAD_POLY[1023-32* 10 -20])^(c[21]&AHEAD_POLY[1023-32* 10 -21])^(c[22]&AHEAD_POLY[1023-32* 10 -22])^(c[23]&AHEAD_POLY[1023-32* 10 -23])^(c[24]&AHEAD_POLY[1023-32* 10 -24])^(c[25]&AHEAD_POLY[1023-32* 10 -25])^(c[26]&AHEAD_POLY[1023-32* 10 -26])^(c[27]&AHEAD_POLY[1023-32* 10 -27])^(c[28]&AHEAD_POLY[1023-32* 10 -28])^(c[29]&AHEAD_POLY[1023-32* 10 -29])^(c[30]&AHEAD_POLY[1023-32* 10 -30])^(c[31]&AHEAD_POLY[1023-32* 10 -31]);
  //   newcrc[11]  = (c[0]&AHEAD_POLY[1023-32* 11 ])^(c[1]&AHEAD_POLY[1023-32* 11 -1])^(c[2]&AHEAD_POLY[1023-32* -2 ])^(c[3]&AHEAD_POLY[1023-32* 11 -3])^(c[4]&AHEAD_POLY[1023-32* 11 -4])^(c[5]&AHEAD_POLY[1023-32* 11 -5])^(c[6]&AHEAD_POLY[1023-32* 11 -6])^(c[7]&AHEAD_POLY[1023-32* 11 -7])^(c[8]&AHEAD_POLY[1023-32* 11 -8])^(c[9]&AHEAD_POLY[1023-32* 11 -9])^(c[10]&AHEAD_POLY[1023-32* 11 -10])^(c[11]&AHEAD_POLY[1023-32* 11 -11])^(c[12]&AHEAD_POLY[1023-32* 11 -12])^(c[13]&AHEAD_POLY[1023-32* 11 -13])^(c[14]&AHEAD_POLY[1023-32* 11 -14])^(c[15]&AHEAD_POLY[1023-32* 11 -15])^(c[16]&AHEAD_POLY[1023-32* 11 -16])^(c[17]&AHEAD_POLY[1023-32* 11 -17])^(c[18]&AHEAD_POLY[1023-32* 11 -18])^(c[19]&AHEAD_POLY[1023-32* 11 -19])^(c[20]&AHEAD_POLY[1023-32* 11 -20])^(c[21]&AHEAD_POLY[1023-32* 11 -21])^(c[22]&AHEAD_POLY[1023-32* 11 -22])^(c[23]&AHEAD_POLY[1023-32* 11 -23])^(c[24]&AHEAD_POLY[1023-32* 11 -24])^(c[25]&AHEAD_POLY[1023-32* 11 -25])^(c[26]&AHEAD_POLY[1023-32* 11 -26])^(c[27]&AHEAD_POLY[1023-32* 11 -27])^(c[28]&AHEAD_POLY[1023-32* 11 -28])^(c[29]&AHEAD_POLY[1023-32* 11 -29])^(c[30]&AHEAD_POLY[1023-32* 11 -30])^(c[31]&AHEAD_POLY[1023-32* 11 -31]);
  //   newcrc[12]  = (c[0]&AHEAD_POLY[1023-32* 12 ])^(c[1]&AHEAD_POLY[1023-32* 12 -1])^(c[2]&AHEAD_POLY[1023-32* -2 ])^(c[3]&AHEAD_POLY[1023-32* 12 -3])^(c[4]&AHEAD_POLY[1023-32* 12 -4])^(c[5]&AHEAD_POLY[1023-32* 12 -5])^(c[6]&AHEAD_POLY[1023-32* 12 -6])^(c[7]&AHEAD_POLY[1023-32* 12 -7])^(c[8]&AHEAD_POLY[1023-32* 12 -8])^(c[9]&AHEAD_POLY[1023-32* 12 -9])^(c[10]&AHEAD_POLY[1023-32* 12 -10])^(c[11]&AHEAD_POLY[1023-32* 12 -11])^(c[12]&AHEAD_POLY[1023-32* 12 -12])^(c[13]&AHEAD_POLY[1023-32* 12 -13])^(c[14]&AHEAD_POLY[1023-32* 12 -14])^(c[15]&AHEAD_POLY[1023-32* 12 -15])^(c[16]&AHEAD_POLY[1023-32* 12 -16])^(c[17]&AHEAD_POLY[1023-32* 12 -17])^(c[18]&AHEAD_POLY[1023-32* 12 -18])^(c[19]&AHEAD_POLY[1023-32* 12 -19])^(c[20]&AHEAD_POLY[1023-32* 12 -20])^(c[21]&AHEAD_POLY[1023-32* 12 -21])^(c[22]&AHEAD_POLY[1023-32* 12 -22])^(c[23]&AHEAD_POLY[1023-32* 12 -23])^(c[24]&AHEAD_POLY[1023-32* 12 -24])^(c[25]&AHEAD_POLY[1023-32* 12 -25])^(c[26]&AHEAD_POLY[1023-32* 12 -26])^(c[27]&AHEAD_POLY[1023-32* 12 -27])^(c[28]&AHEAD_POLY[1023-32* 12 -28])^(c[29]&AHEAD_POLY[1023-32* 12 -29])^(c[30]&AHEAD_POLY[1023-32* 12 -30])^(c[31]&AHEAD_POLY[1023-32* 12 -31]);
  //   newcrc[13]  = (c[0]&AHEAD_POLY[1023-32* 13 ])^(c[1]&AHEAD_POLY[1023-32* 13 -1])^(c[2]&AHEAD_POLY[1023-32* -2 ])^(c[3]&AHEAD_POLY[1023-32* 13 -3])^(c[4]&AHEAD_POLY[1023-32* 13 -4])^(c[5]&AHEAD_POLY[1023-32* 13 -5])^(c[6]&AHEAD_POLY[1023-32* 13 -6])^(c[7]&AHEAD_POLY[1023-32* 13 -7])^(c[8]&AHEAD_POLY[1023-32* 13 -8])^(c[9]&AHEAD_POLY[1023-32* 13 -9])^(c[10]&AHEAD_POLY[1023-32* 13 -10])^(c[11]&AHEAD_POLY[1023-32* 13 -11])^(c[12]&AHEAD_POLY[1023-32* 13 -12])^(c[13]&AHEAD_POLY[1023-32* 13 -13])^(c[14]&AHEAD_POLY[1023-32* 13 -14])^(c[15]&AHEAD_POLY[1023-32* 13 -15])^(c[16]&AHEAD_POLY[1023-32* 13 -16])^(c[17]&AHEAD_POLY[1023-32* 13 -17])^(c[18]&AHEAD_POLY[1023-32* 13 -18])^(c[19]&AHEAD_POLY[1023-32* 13 -19])^(c[20]&AHEAD_POLY[1023-32* 13 -20])^(c[21]&AHEAD_POLY[1023-32* 13 -21])^(c[22]&AHEAD_POLY[1023-32* 13 -22])^(c[23]&AHEAD_POLY[1023-32* 13 -23])^(c[24]&AHEAD_POLY[1023-32* 13 -24])^(c[25]&AHEAD_POLY[1023-32* 13 -25])^(c[26]&AHEAD_POLY[1023-32* 13 -26])^(c[27]&AHEAD_POLY[1023-32* 13 -27])^(c[28]&AHEAD_POLY[1023-32* 13 -28])^(c[29]&AHEAD_POLY[1023-32* 13 -29])^(c[30]&AHEAD_POLY[1023-32* 13 -30])^(c[31]&AHEAD_POLY[1023-32* 13 -31]);
  //   newcrc[14]  = (c[0]&AHEAD_POLY[1023-32* 14 ])^(c[1]&AHEAD_POLY[1023-32* 14 -1])^(c[2]&AHEAD_POLY[1023-32* -2 ])^(c[3]&AHEAD_POLY[1023-32* 14 -3])^(c[4]&AHEAD_POLY[1023-32* 14 -4])^(c[5]&AHEAD_POLY[1023-32* 14 -5])^(c[6]&AHEAD_POLY[1023-32* 14 -6])^(c[7]&AHEAD_POLY[1023-32* 14 -7])^(c[8]&AHEAD_POLY[1023-32* 14 -8])^(c[9]&AHEAD_POLY[1023-32* 14 -9])^(c[10]&AHEAD_POLY[1023-32* 14 -10])^(c[11]&AHEAD_POLY[1023-32* 14 -11])^(c[12]&AHEAD_POLY[1023-32* 14 -12])^(c[13]&AHEAD_POLY[1023-32* 14 -13])^(c[14]&AHEAD_POLY[1023-32* 14 -14])^(c[15]&AHEAD_POLY[1023-32* 14 -15])^(c[16]&AHEAD_POLY[1023-32* 14 -16])^(c[17]&AHEAD_POLY[1023-32* 14 -17])^(c[18]&AHEAD_POLY[1023-32* 14 -18])^(c[19]&AHEAD_POLY[1023-32* 14 -19])^(c[20]&AHEAD_POLY[1023-32* 14 -20])^(c[21]&AHEAD_POLY[1023-32* 14 -21])^(c[22]&AHEAD_POLY[1023-32* 14 -22])^(c[23]&AHEAD_POLY[1023-32* 14 -23])^(c[24]&AHEAD_POLY[1023-32* 14 -24])^(c[25]&AHEAD_POLY[1023-32* 14 -25])^(c[26]&AHEAD_POLY[1023-32* 14 -26])^(c[27]&AHEAD_POLY[1023-32* 14 -27])^(c[28]&AHEAD_POLY[1023-32* 14 -28])^(c[29]&AHEAD_POLY[1023-32* 14 -29])^(c[30]&AHEAD_POLY[1023-32* 14 -30])^(c[31]&AHEAD_POLY[1023-32* 14 -31]);
  //   newcrc[15]  = (c[0]&AHEAD_POLY[1023-32* 15 ])^(c[1]&AHEAD_POLY[1023-32* 15 -1])^(c[2]&AHEAD_POLY[1023-32* -2 ])^(c[3]&AHEAD_POLY[1023-32* 15 -3])^(c[4]&AHEAD_POLY[1023-32* 15 -4])^(c[5]&AHEAD_POLY[1023-32* 15 -5])^(c[6]&AHEAD_POLY[1023-32* 15 -6])^(c[7]&AHEAD_POLY[1023-32* 15 -7])^(c[8]&AHEAD_POLY[1023-32* 15 -8])^(c[9]&AHEAD_POLY[1023-32* 15 -9])^(c[10]&AHEAD_POLY[1023-32* 15 -10])^(c[11]&AHEAD_POLY[1023-32* 15 -11])^(c[12]&AHEAD_POLY[1023-32* 15 -12])^(c[13]&AHEAD_POLY[1023-32* 15 -13])^(c[14]&AHEAD_POLY[1023-32* 15 -14])^(c[15]&AHEAD_POLY[1023-32* 15 -15])^(c[16]&AHEAD_POLY[1023-32* 15 -16])^(c[17]&AHEAD_POLY[1023-32* 15 -17])^(c[18]&AHEAD_POLY[1023-32* 15 -18])^(c[19]&AHEAD_POLY[1023-32* 15 -19])^(c[20]&AHEAD_POLY[1023-32* 15 -20])^(c[21]&AHEAD_POLY[1023-32* 15 -21])^(c[22]&AHEAD_POLY[1023-32* 15 -22])^(c[23]&AHEAD_POLY[1023-32* 15 -23])^(c[24]&AHEAD_POLY[1023-32* 15 -24])^(c[25]&AHEAD_POLY[1023-32* 15 -25])^(c[26]&AHEAD_POLY[1023-32* 15 -26])^(c[27]&AHEAD_POLY[1023-32* 15 -27])^(c[28]&AHEAD_POLY[1023-32* 15 -28])^(c[29]&AHEAD_POLY[1023-32* 15 -29])^(c[30]&AHEAD_POLY[1023-32* 15 -30])^(c[31]&AHEAD_POLY[1023-32* 15 -31]);
  //   newcrc[16]  = (c[0]&AHEAD_POLY[1023-32* 16 ])^(c[1]&AHEAD_POLY[1023-32* 16 -1])^(c[2]&AHEAD_POLY[1023-32* -2 ])^(c[3]&AHEAD_POLY[1023-32* 16 -3])^(c[4]&AHEAD_POLY[1023-32* 16 -4])^(c[5]&AHEAD_POLY[1023-32* 16 -5])^(c[6]&AHEAD_POLY[1023-32* 16 -6])^(c[7]&AHEAD_POLY[1023-32* 16 -7])^(c[8]&AHEAD_POLY[1023-32* 16 -8])^(c[9]&AHEAD_POLY[1023-32* 16 -9])^(c[10]&AHEAD_POLY[1023-32* 16 -10])^(c[11]&AHEAD_POLY[1023-32* 16 -11])^(c[12]&AHEAD_POLY[1023-32* 16 -12])^(c[13]&AHEAD_POLY[1023-32* 16 -13])^(c[14]&AHEAD_POLY[1023-32* 16 -14])^(c[15]&AHEAD_POLY[1023-32* 16 -15])^(c[16]&AHEAD_POLY[1023-32* 16 -16])^(c[17]&AHEAD_POLY[1023-32* 16 -17])^(c[18]&AHEAD_POLY[1023-32* 16 -18])^(c[19]&AHEAD_POLY[1023-32* 16 -19])^(c[20]&AHEAD_POLY[1023-32* 16 -20])^(c[21]&AHEAD_POLY[1023-32* 16 -21])^(c[22]&AHEAD_POLY[1023-32* 16 -22])^(c[23]&AHEAD_POLY[1023-32* 16 -23])^(c[24]&AHEAD_POLY[1023-32* 16 -24])^(c[25]&AHEAD_POLY[1023-32* 16 -25])^(c[26]&AHEAD_POLY[1023-32* 16 -26])^(c[27]&AHEAD_POLY[1023-32* 16 -27])^(c[28]&AHEAD_POLY[1023-32* 16 -28])^(c[29]&AHEAD_POLY[1023-32* 16 -29])^(c[30]&AHEAD_POLY[1023-32* 16 -30])^(c[31]&AHEAD_POLY[1023-32* 16 -31]);
  //   newcrc[17]  = (c[0]&AHEAD_POLY[1023-32* 17 ])^(c[1]&AHEAD_POLY[1023-32* 17 -1])^(c[2]&AHEAD_POLY[1023-32* -2 ])^(c[3]&AHEAD_POLY[1023-32* 17 -3])^(c[4]&AHEAD_POLY[1023-32* 17 -4])^(c[5]&AHEAD_POLY[1023-32* 17 -5])^(c[6]&AHEAD_POLY[1023-32* 17 -6])^(c[7]&AHEAD_POLY[1023-32* 17 -7])^(c[8]&AHEAD_POLY[1023-32* 17 -8])^(c[9]&AHEAD_POLY[1023-32* 17 -9])^(c[10]&AHEAD_POLY[1023-32* 17 -10])^(c[11]&AHEAD_POLY[1023-32* 17 -11])^(c[12]&AHEAD_POLY[1023-32* 17 -12])^(c[13]&AHEAD_POLY[1023-32* 17 -13])^(c[14]&AHEAD_POLY[1023-32* 17 -14])^(c[15]&AHEAD_POLY[1023-32* 17 -15])^(c[16]&AHEAD_POLY[1023-32* 17 -16])^(c[17]&AHEAD_POLY[1023-32* 17 -17])^(c[18]&AHEAD_POLY[1023-32* 17 -18])^(c[19]&AHEAD_POLY[1023-32* 17 -19])^(c[20]&AHEAD_POLY[1023-32* 17 -20])^(c[21]&AHEAD_POLY[1023-32* 17 -21])^(c[22]&AHEAD_POLY[1023-32* 17 -22])^(c[23]&AHEAD_POLY[1023-32* 17 -23])^(c[24]&AHEAD_POLY[1023-32* 17 -24])^(c[25]&AHEAD_POLY[1023-32* 17 -25])^(c[26]&AHEAD_POLY[1023-32* 17 -26])^(c[27]&AHEAD_POLY[1023-32* 17 -27])^(c[28]&AHEAD_POLY[1023-32* 17 -28])^(c[29]&AHEAD_POLY[1023-32* 17 -29])^(c[30]&AHEAD_POLY[1023-32* 17 -30])^(c[31]&AHEAD_POLY[1023-32* 17 -31]);
  //   newcrc[18]  = (c[0]&AHEAD_POLY[1023-32* 18 ])^(c[1]&AHEAD_POLY[1023-32* 18 -1])^(c[2]&AHEAD_POLY[1023-32* -2 ])^(c[3]&AHEAD_POLY[1023-32* 18 -3])^(c[4]&AHEAD_POLY[1023-32* 18 -4])^(c[5]&AHEAD_POLY[1023-32* 18 -5])^(c[6]&AHEAD_POLY[1023-32* 18 -6])^(c[7]&AHEAD_POLY[1023-32* 18 -7])^(c[8]&AHEAD_POLY[1023-32* 18 -8])^(c[9]&AHEAD_POLY[1023-32* 18 -9])^(c[10]&AHEAD_POLY[1023-32* 18 -10])^(c[11]&AHEAD_POLY[1023-32* 18 -11])^(c[12]&AHEAD_POLY[1023-32* 18 -12])^(c[13]&AHEAD_POLY[1023-32* 18 -13])^(c[14]&AHEAD_POLY[1023-32* 18 -14])^(c[15]&AHEAD_POLY[1023-32* 18 -15])^(c[16]&AHEAD_POLY[1023-32* 18 -16])^(c[17]&AHEAD_POLY[1023-32* 18 -17])^(c[18]&AHEAD_POLY[1023-32* 18 -18])^(c[19]&AHEAD_POLY[1023-32* 18 -19])^(c[20]&AHEAD_POLY[1023-32* 18 -20])^(c[21]&AHEAD_POLY[1023-32* 18 -21])^(c[22]&AHEAD_POLY[1023-32* 18 -22])^(c[23]&AHEAD_POLY[1023-32* 18 -23])^(c[24]&AHEAD_POLY[1023-32* 18 -24])^(c[25]&AHEAD_POLY[1023-32* 18 -25])^(c[26]&AHEAD_POLY[1023-32* 18 -26])^(c[27]&AHEAD_POLY[1023-32* 18 -27])^(c[28]&AHEAD_POLY[1023-32* 18 -28])^(c[29]&AHEAD_POLY[1023-32* 18 -29])^(c[30]&AHEAD_POLY[1023-32* 18 -30])^(c[31]&AHEAD_POLY[1023-32* 18 -31]);
  //   newcrc[19]  = (c[0]&AHEAD_POLY[1023-32* 19 ])^(c[1]&AHEAD_POLY[1023-32* 19 -1])^(c[2]&AHEAD_POLY[1023-32* -2 ])^(c[3]&AHEAD_POLY[1023-32* 19 -3])^(c[4]&AHEAD_POLY[1023-32* 19 -4])^(c[5]&AHEAD_POLY[1023-32* 19 -5])^(c[6]&AHEAD_POLY[1023-32* 19 -6])^(c[7]&AHEAD_POLY[1023-32* 19 -7])^(c[8]&AHEAD_POLY[1023-32* 19 -8])^(c[9]&AHEAD_POLY[1023-32* 19 -9])^(c[10]&AHEAD_POLY[1023-32* 19 -10])^(c[11]&AHEAD_POLY[1023-32* 19 -11])^(c[12]&AHEAD_POLY[1023-32* 19 -12])^(c[13]&AHEAD_POLY[1023-32* 19 -13])^(c[14]&AHEAD_POLY[1023-32* 19 -14])^(c[15]&AHEAD_POLY[1023-32* 19 -15])^(c[16]&AHEAD_POLY[1023-32* 19 -16])^(c[17]&AHEAD_POLY[1023-32* 19 -17])^(c[18]&AHEAD_POLY[1023-32* 19 -18])^(c[19]&AHEAD_POLY[1023-32* 19 -19])^(c[20]&AHEAD_POLY[1023-32* 19 -20])^(c[21]&AHEAD_POLY[1023-32* 19 -21])^(c[22]&AHEAD_POLY[1023-32* 19 -22])^(c[23]&AHEAD_POLY[1023-32* 19 -23])^(c[24]&AHEAD_POLY[1023-32* 19 -24])^(c[25]&AHEAD_POLY[1023-32* 19 -25])^(c[26]&AHEAD_POLY[1023-32* 19 -26])^(c[27]&AHEAD_POLY[1023-32* 19 -27])^(c[28]&AHEAD_POLY[1023-32* 19 -28])^(c[29]&AHEAD_POLY[1023-32* 19 -29])^(c[30]&AHEAD_POLY[1023-32* 19 -30])^(c[31]&AHEAD_POLY[1023-32* 19 -31]);
  //   newcrc[20]  = (c[0]&AHEAD_POLY[1023-32* 20 ])^(c[1]&AHEAD_POLY[1023-32* 20 -1])^(c[2]&AHEAD_POLY[1023-32* -2 ])^(c[3]&AHEAD_POLY[1023-32* 20 -3])^(c[4]&AHEAD_POLY[1023-32* 20 -4])^(c[5]&AHEAD_POLY[1023-32* 20 -5])^(c[6]&AHEAD_POLY[1023-32* 20 -6])^(c[7]&AHEAD_POLY[1023-32* 20 -7])^(c[8]&AHEAD_POLY[1023-32* 20 -8])^(c[9]&AHEAD_POLY[1023-32* 20 -9])^(c[10]&AHEAD_POLY[1023-32* 20 -10])^(c[11]&AHEAD_POLY[1023-32* 20 -11])^(c[12]&AHEAD_POLY[1023-32* 20 -12])^(c[13]&AHEAD_POLY[1023-32* 20 -13])^(c[14]&AHEAD_POLY[1023-32* 20 -14])^(c[15]&AHEAD_POLY[1023-32* 20 -15])^(c[16]&AHEAD_POLY[1023-32* 20 -16])^(c[17]&AHEAD_POLY[1023-32* 20 -17])^(c[18]&AHEAD_POLY[1023-32* 20 -18])^(c[19]&AHEAD_POLY[1023-32* 20 -19])^(c[20]&AHEAD_POLY[1023-32* 20 -20])^(c[21]&AHEAD_POLY[1023-32* 20 -21])^(c[22]&AHEAD_POLY[1023-32* 20 -22])^(c[23]&AHEAD_POLY[1023-32* 20 -23])^(c[24]&AHEAD_POLY[1023-32* 20 -24])^(c[25]&AHEAD_POLY[1023-32* 20 -25])^(c[26]&AHEAD_POLY[1023-32* 20 -26])^(c[27]&AHEAD_POLY[1023-32* 20 -27])^(c[28]&AHEAD_POLY[1023-32* 20 -28])^(c[29]&AHEAD_POLY[1023-32* 20 -29])^(c[30]&AHEAD_POLY[1023-32* 20 -30])^(c[31]&AHEAD_POLY[1023-32* 20 -31]);
  //   newcrc[21]  = (c[0]&AHEAD_POLY[1023-32* 21 ])^(c[1]&AHEAD_POLY[1023-32* 21 -1])^(c[2]&AHEAD_POLY[1023-32* -2 ])^(c[3]&AHEAD_POLY[1023-32* 21 -3])^(c[4]&AHEAD_POLY[1023-32* 21 -4])^(c[5]&AHEAD_POLY[1023-32* 21 -5])^(c[6]&AHEAD_POLY[1023-32* 21 -6])^(c[7]&AHEAD_POLY[1023-32* 21 -7])^(c[8]&AHEAD_POLY[1023-32* 21 -8])^(c[9]&AHEAD_POLY[1023-32* 21 -9])^(c[10]&AHEAD_POLY[1023-32* 21 -10])^(c[11]&AHEAD_POLY[1023-32* 21 -11])^(c[12]&AHEAD_POLY[1023-32* 21 -12])^(c[13]&AHEAD_POLY[1023-32* 21 -13])^(c[14]&AHEAD_POLY[1023-32* 21 -14])^(c[15]&AHEAD_POLY[1023-32* 21 -15])^(c[16]&AHEAD_POLY[1023-32* 21 -16])^(c[17]&AHEAD_POLY[1023-32* 21 -17])^(c[18]&AHEAD_POLY[1023-32* 21 -18])^(c[19]&AHEAD_POLY[1023-32* 21 -19])^(c[20]&AHEAD_POLY[1023-32* 21 -20])^(c[21]&AHEAD_POLY[1023-32* 21 -21])^(c[22]&AHEAD_POLY[1023-32* 21 -22])^(c[23]&AHEAD_POLY[1023-32* 21 -23])^(c[24]&AHEAD_POLY[1023-32* 21 -24])^(c[25]&AHEAD_POLY[1023-32* 21 -25])^(c[26]&AHEAD_POLY[1023-32* 21 -26])^(c[27]&AHEAD_POLY[1023-32* 21 -27])^(c[28]&AHEAD_POLY[1023-32* 21 -28])^(c[29]&AHEAD_POLY[1023-32* 21 -29])^(c[30]&AHEAD_POLY[1023-32* 21 -30])^(c[31]&AHEAD_POLY[1023-32* 21 -31]);
  //   newcrc[22]  = (c[0]&AHEAD_POLY[1023-32* 22 ])^(c[1]&AHEAD_POLY[1023-32* 22 -1])^(c[2]&AHEAD_POLY[1023-32* -2 ])^(c[3]&AHEAD_POLY[1023-32* 22 -3])^(c[4]&AHEAD_POLY[1023-32* 22 -4])^(c[5]&AHEAD_POLY[1023-32* 22 -5])^(c[6]&AHEAD_POLY[1023-32* 22 -6])^(c[7]&AHEAD_POLY[1023-32* 22 -7])^(c[8]&AHEAD_POLY[1023-32* 22 -8])^(c[9]&AHEAD_POLY[1023-32* 22 -9])^(c[10]&AHEAD_POLY[1023-32* 22 -10])^(c[11]&AHEAD_POLY[1023-32* 22 -11])^(c[12]&AHEAD_POLY[1023-32* 22 -12])^(c[13]&AHEAD_POLY[1023-32* 22 -13])^(c[14]&AHEAD_POLY[1023-32* 22 -14])^(c[15]&AHEAD_POLY[1023-32* 22 -15])^(c[16]&AHEAD_POLY[1023-32* 22 -16])^(c[17]&AHEAD_POLY[1023-32* 22 -17])^(c[18]&AHEAD_POLY[1023-32* 22 -18])^(c[19]&AHEAD_POLY[1023-32* 22 -19])^(c[20]&AHEAD_POLY[1023-32* 22 -20])^(c[21]&AHEAD_POLY[1023-32* 22 -21])^(c[22]&AHEAD_POLY[1023-32* 22 -22])^(c[23]&AHEAD_POLY[1023-32* 22 -23])^(c[24]&AHEAD_POLY[1023-32* 22 -24])^(c[25]&AHEAD_POLY[1023-32* 22 -25])^(c[26]&AHEAD_POLY[1023-32* 22 -26])^(c[27]&AHEAD_POLY[1023-32* 22 -27])^(c[28]&AHEAD_POLY[1023-32* 22 -28])^(c[29]&AHEAD_POLY[1023-32* 22 -29])^(c[30]&AHEAD_POLY[1023-32* 22 -30])^(c[31]&AHEAD_POLY[1023-32* 22 -31]);
  //   newcrc[23]  = (c[0]&AHEAD_POLY[1023-32* 23 ])^(c[1]&AHEAD_POLY[1023-32* 23 -1])^(c[2]&AHEAD_POLY[1023-32* -2 ])^(c[3]&AHEAD_POLY[1023-32* 23 -3])^(c[4]&AHEAD_POLY[1023-32* 23 -4])^(c[5]&AHEAD_POLY[1023-32* 23 -5])^(c[6]&AHEAD_POLY[1023-32* 23 -6])^(c[7]&AHEAD_POLY[1023-32* 23 -7])^(c[8]&AHEAD_POLY[1023-32* 23 -8])^(c[9]&AHEAD_POLY[1023-32* 23 -9])^(c[10]&AHEAD_POLY[1023-32* 23 -10])^(c[11]&AHEAD_POLY[1023-32* 23 -11])^(c[12]&AHEAD_POLY[1023-32* 23 -12])^(c[13]&AHEAD_POLY[1023-32* 23 -13])^(c[14]&AHEAD_POLY[1023-32* 23 -14])^(c[15]&AHEAD_POLY[1023-32* 23 -15])^(c[16]&AHEAD_POLY[1023-32* 23 -16])^(c[17]&AHEAD_POLY[1023-32* 23 -17])^(c[18]&AHEAD_POLY[1023-32* 23 -18])^(c[19]&AHEAD_POLY[1023-32* 23 -19])^(c[20]&AHEAD_POLY[1023-32* 23 -20])^(c[21]&AHEAD_POLY[1023-32* 23 -21])^(c[22]&AHEAD_POLY[1023-32* 23 -22])^(c[23]&AHEAD_POLY[1023-32* 23 -23])^(c[24]&AHEAD_POLY[1023-32* 23 -24])^(c[25]&AHEAD_POLY[1023-32* 23 -25])^(c[26]&AHEAD_POLY[1023-32* 23 -26])^(c[27]&AHEAD_POLY[1023-32* 23 -27])^(c[28]&AHEAD_POLY[1023-32* 23 -28])^(c[29]&AHEAD_POLY[1023-32* 23 -29])^(c[30]&AHEAD_POLY[1023-32* 23 -30])^(c[31]&AHEAD_POLY[1023-32* 23 -31]);
  //   newcrc[24]  = (c[0]&AHEAD_POLY[1023-32* 24 ])^(c[1]&AHEAD_POLY[1023-32* 24 -1])^(c[2]&AHEAD_POLY[1023-32* -2 ])^(c[3]&AHEAD_POLY[1023-32* 24 -3])^(c[4]&AHEAD_POLY[1023-32* 24 -4])^(c[5]&AHEAD_POLY[1023-32* 24 -5])^(c[6]&AHEAD_POLY[1023-32* 24 -6])^(c[7]&AHEAD_POLY[1023-32* 24 -7])^(c[8]&AHEAD_POLY[1023-32* 24 -8])^(c[9]&AHEAD_POLY[1023-32* 24 -9])^(c[10]&AHEAD_POLY[1023-32* 24 -10])^(c[11]&AHEAD_POLY[1023-32* 24 -11])^(c[12]&AHEAD_POLY[1023-32* 24 -12])^(c[13]&AHEAD_POLY[1023-32* 24 -13])^(c[14]&AHEAD_POLY[1023-32* 24 -14])^(c[15]&AHEAD_POLY[1023-32* 24 -15])^(c[16]&AHEAD_POLY[1023-32* 24 -16])^(c[17]&AHEAD_POLY[1023-32* 24 -17])^(c[18]&AHEAD_POLY[1023-32* 24 -18])^(c[19]&AHEAD_POLY[1023-32* 24 -19])^(c[20]&AHEAD_POLY[1023-32* 24 -20])^(c[21]&AHEAD_POLY[1023-32* 24 -21])^(c[22]&AHEAD_POLY[1023-32* 24 -22])^(c[23]&AHEAD_POLY[1023-32* 24 -23])^(c[24]&AHEAD_POLY[1023-32* 24 -24])^(c[25]&AHEAD_POLY[1023-32* 24 -25])^(c[26]&AHEAD_POLY[1023-32* 24 -26])^(c[27]&AHEAD_POLY[1023-32* 24 -27])^(c[28]&AHEAD_POLY[1023-32* 24 -28])^(c[29]&AHEAD_POLY[1023-32* 24 -29])^(c[30]&AHEAD_POLY[1023-32* 24 -30])^(c[31]&AHEAD_POLY[1023-32* 24 -31]);
  //   newcrc[25]  = (c[0]&AHEAD_POLY[1023-32* 25 ])^(c[1]&AHEAD_POLY[1023-32* 25 -1])^(c[2]&AHEAD_POLY[1023-32* -2 ])^(c[3]&AHEAD_POLY[1023-32* 25 -3])^(c[4]&AHEAD_POLY[1023-32* 25 -4])^(c[5]&AHEAD_POLY[1023-32* 25 -5])^(c[6]&AHEAD_POLY[1023-32* 25 -6])^(c[7]&AHEAD_POLY[1023-32* 25 -7])^(c[8]&AHEAD_POLY[1023-32* 25 -8])^(c[9]&AHEAD_POLY[1023-32* 25 -9])^(c[10]&AHEAD_POLY[1023-32* 25 -10])^(c[11]&AHEAD_POLY[1023-32* 25 -11])^(c[12]&AHEAD_POLY[1023-32* 25 -12])^(c[13]&AHEAD_POLY[1023-32* 25 -13])^(c[14]&AHEAD_POLY[1023-32* 25 -14])^(c[15]&AHEAD_POLY[1023-32* 25 -15])^(c[16]&AHEAD_POLY[1023-32* 25 -16])^(c[17]&AHEAD_POLY[1023-32* 25 -17])^(c[18]&AHEAD_POLY[1023-32* 25 -18])^(c[19]&AHEAD_POLY[1023-32* 25 -19])^(c[20]&AHEAD_POLY[1023-32* 25 -20])^(c[21]&AHEAD_POLY[1023-32* 25 -21])^(c[22]&AHEAD_POLY[1023-32* 25 -22])^(c[23]&AHEAD_POLY[1023-32* 25 -23])^(c[24]&AHEAD_POLY[1023-32* 25 -24])^(c[25]&AHEAD_POLY[1023-32* 25 -25])^(c[26]&AHEAD_POLY[1023-32* 25 -26])^(c[27]&AHEAD_POLY[1023-32* 25 -27])^(c[28]&AHEAD_POLY[1023-32* 25 -28])^(c[29]&AHEAD_POLY[1023-32* 25 -29])^(c[30]&AHEAD_POLY[1023-32* 25 -30])^(c[31]&AHEAD_POLY[1023-32* 25 -31]);
  //   newcrc[26]  = (c[0]&AHEAD_POLY[1023-32* 26 ])^(c[1]&AHEAD_POLY[1023-32* 26 -1])^(c[2]&AHEAD_POLY[1023-32* -2 ])^(c[3]&AHEAD_POLY[1023-32* 26 -3])^(c[4]&AHEAD_POLY[1023-32* 26 -4])^(c[5]&AHEAD_POLY[1023-32* 26 -5])^(c[6]&AHEAD_POLY[1023-32* 26 -6])^(c[7]&AHEAD_POLY[1023-32* 26 -7])^(c[8]&AHEAD_POLY[1023-32* 26 -8])^(c[9]&AHEAD_POLY[1023-32* 26 -9])^(c[10]&AHEAD_POLY[1023-32* 26 -10])^(c[11]&AHEAD_POLY[1023-32* 26 -11])^(c[12]&AHEAD_POLY[1023-32* 26 -12])^(c[13]&AHEAD_POLY[1023-32* 26 -13])^(c[14]&AHEAD_POLY[1023-32* 26 -14])^(c[15]&AHEAD_POLY[1023-32* 26 -15])^(c[16]&AHEAD_POLY[1023-32* 26 -16])^(c[17]&AHEAD_POLY[1023-32* 26 -17])^(c[18]&AHEAD_POLY[1023-32* 26 -18])^(c[19]&AHEAD_POLY[1023-32* 26 -19])^(c[20]&AHEAD_POLY[1023-32* 26 -20])^(c[21]&AHEAD_POLY[1023-32* 26 -21])^(c[22]&AHEAD_POLY[1023-32* 26 -22])^(c[23]&AHEAD_POLY[1023-32* 26 -23])^(c[24]&AHEAD_POLY[1023-32* 26 -24])^(c[25]&AHEAD_POLY[1023-32* 26 -25])^(c[26]&AHEAD_POLY[1023-32* 26 -26])^(c[27]&AHEAD_POLY[1023-32* 26 -27])^(c[28]&AHEAD_POLY[1023-32* 26 -28])^(c[29]&AHEAD_POLY[1023-32* 26 -29])^(c[30]&AHEAD_POLY[1023-32* 26 -30])^(c[31]&AHEAD_POLY[1023-32* 26 -31]);
  //   newcrc[27]  = (c[0]&AHEAD_POLY[1023-32* 27 ])^(c[1]&AHEAD_POLY[1023-32* 27 -1])^(c[2]&AHEAD_POLY[1023-32* -2 ])^(c[3]&AHEAD_POLY[1023-32* 27 -3])^(c[4]&AHEAD_POLY[1023-32* 27 -4])^(c[5]&AHEAD_POLY[1023-32* 27 -5])^(c[6]&AHEAD_POLY[1023-32* 27 -6])^(c[7]&AHEAD_POLY[1023-32* 27 -7])^(c[8]&AHEAD_POLY[1023-32* 27 -8])^(c[9]&AHEAD_POLY[1023-32* 27 -9])^(c[10]&AHEAD_POLY[1023-32* 27 -10])^(c[11]&AHEAD_POLY[1023-32* 27 -11])^(c[12]&AHEAD_POLY[1023-32* 27 -12])^(c[13]&AHEAD_POLY[1023-32* 27 -13])^(c[14]&AHEAD_POLY[1023-32* 27 -14])^(c[15]&AHEAD_POLY[1023-32* 27 -15])^(c[16]&AHEAD_POLY[1023-32* 27 -16])^(c[17]&AHEAD_POLY[1023-32* 27 -17])^(c[18]&AHEAD_POLY[1023-32* 27 -18])^(c[19]&AHEAD_POLY[1023-32* 27 -19])^(c[20]&AHEAD_POLY[1023-32* 27 -20])^(c[21]&AHEAD_POLY[1023-32* 27 -21])^(c[22]&AHEAD_POLY[1023-32* 27 -22])^(c[23]&AHEAD_POLY[1023-32* 27 -23])^(c[24]&AHEAD_POLY[1023-32* 27 -24])^(c[25]&AHEAD_POLY[1023-32* 27 -25])^(c[26]&AHEAD_POLY[1023-32* 27 -26])^(c[27]&AHEAD_POLY[1023-32* 27 -27])^(c[28]&AHEAD_POLY[1023-32* 27 -28])^(c[29]&AHEAD_POLY[1023-32* 27 -29])^(c[30]&AHEAD_POLY[1023-32* 27 -30])^(c[31]&AHEAD_POLY[1023-32* 27 -31]);
  //   newcrc[28]  = (c[0]&AHEAD_POLY[1023-32* 28 ])^(c[1]&AHEAD_POLY[1023-32* 28 -1])^(c[2]&AHEAD_POLY[1023-32* -2 ])^(c[3]&AHEAD_POLY[1023-32* 28 -3])^(c[4]&AHEAD_POLY[1023-32* 28 -4])^(c[5]&AHEAD_POLY[1023-32* 28 -5])^(c[6]&AHEAD_POLY[1023-32* 28 -6])^(c[7]&AHEAD_POLY[1023-32* 28 -7])^(c[8]&AHEAD_POLY[1023-32* 28 -8])^(c[9]&AHEAD_POLY[1023-32* 28 -9])^(c[10]&AHEAD_POLY[1023-32* 28 -10])^(c[11]&AHEAD_POLY[1023-32* 28 -11])^(c[12]&AHEAD_POLY[1023-32* 28 -12])^(c[13]&AHEAD_POLY[1023-32* 28 -13])^(c[14]&AHEAD_POLY[1023-32* 28 -14])^(c[15]&AHEAD_POLY[1023-32* 28 -15])^(c[16]&AHEAD_POLY[1023-32* 28 -16])^(c[17]&AHEAD_POLY[1023-32* 28 -17])^(c[18]&AHEAD_POLY[1023-32* 28 -18])^(c[19]&AHEAD_POLY[1023-32* 28 -19])^(c[20]&AHEAD_POLY[1023-32* 28 -20])^(c[21]&AHEAD_POLY[1023-32* 28 -21])^(c[22]&AHEAD_POLY[1023-32* 28 -22])^(c[23]&AHEAD_POLY[1023-32* 28 -23])^(c[24]&AHEAD_POLY[1023-32* 28 -24])^(c[25]&AHEAD_POLY[1023-32* 28 -25])^(c[26]&AHEAD_POLY[1023-32* 28 -26])^(c[27]&AHEAD_POLY[1023-32* 28 -27])^(c[28]&AHEAD_POLY[1023-32* 28 -28])^(c[29]&AHEAD_POLY[1023-32* 28 -29])^(c[30]&AHEAD_POLY[1023-32* 28 -30])^(c[31]&AHEAD_POLY[1023-32* 28 -31]);
  //   newcrc[29]  = (c[0]&AHEAD_POLY[1023-32* 29 ])^(c[1]&AHEAD_POLY[1023-32* 29 -1])^(c[2]&AHEAD_POLY[1023-32* -2 ])^(c[3]&AHEAD_POLY[1023-32* 29 -3])^(c[4]&AHEAD_POLY[1023-32* 29 -4])^(c[5]&AHEAD_POLY[1023-32* 29 -5])^(c[6]&AHEAD_POLY[1023-32* 29 -6])^(c[7]&AHEAD_POLY[1023-32* 29 -7])^(c[8]&AHEAD_POLY[1023-32* 29 -8])^(c[9]&AHEAD_POLY[1023-32* 29 -9])^(c[10]&AHEAD_POLY[1023-32* 29 -10])^(c[11]&AHEAD_POLY[1023-32* 29 -11])^(c[12]&AHEAD_POLY[1023-32* 29 -12])^(c[13]&AHEAD_POLY[1023-32* 29 -13])^(c[14]&AHEAD_POLY[1023-32* 29 -14])^(c[15]&AHEAD_POLY[1023-32* 29 -15])^(c[16]&AHEAD_POLY[1023-32* 29 -16])^(c[17]&AHEAD_POLY[1023-32* 29 -17])^(c[18]&AHEAD_POLY[1023-32* 29 -18])^(c[19]&AHEAD_POLY[1023-32* 29 -19])^(c[20]&AHEAD_POLY[1023-32* 29 -20])^(c[21]&AHEAD_POLY[1023-32* 29 -21])^(c[22]&AHEAD_POLY[1023-32* 29 -22])^(c[23]&AHEAD_POLY[1023-32* 29 -23])^(c[24]&AHEAD_POLY[1023-32* 29 -24])^(c[25]&AHEAD_POLY[1023-32* 29 -25])^(c[26]&AHEAD_POLY[1023-32* 29 -26])^(c[27]&AHEAD_POLY[1023-32* 29 -27])^(c[28]&AHEAD_POLY[1023-32* 29 -28])^(c[29]&AHEAD_POLY[1023-32* 29 -29])^(c[30]&AHEAD_POLY[1023-32* 29 -30])^(c[31]&AHEAD_POLY[1023-32* 29 -31]);
  //   newcrc[30]  = (c[0]&AHEAD_POLY[1023-32* 30 ])^(c[1]&AHEAD_POLY[1023-32* 30 -1])^(c[2]&AHEAD_POLY[1023-32* -2 ])^(c[3]&AHEAD_POLY[1023-32* 30 -3])^(c[4]&AHEAD_POLY[1023-32* 30 -4])^(c[5]&AHEAD_POLY[1023-32* 30 -5])^(c[6]&AHEAD_POLY[1023-32* 30 -6])^(c[7]&AHEAD_POLY[1023-32* 30 -7])^(c[8]&AHEAD_POLY[1023-32* 30 -8])^(c[9]&AHEAD_POLY[1023-32* 30 -9])^(c[10]&AHEAD_POLY[1023-32* 30 -10])^(c[11]&AHEAD_POLY[1023-32* 30 -11])^(c[12]&AHEAD_POLY[1023-32* 30 -12])^(c[13]&AHEAD_POLY[1023-32* 30 -13])^(c[14]&AHEAD_POLY[1023-32* 30 -14])^(c[15]&AHEAD_POLY[1023-32* 30 -15])^(c[16]&AHEAD_POLY[1023-32* 30 -16])^(c[17]&AHEAD_POLY[1023-32* 30 -17])^(c[18]&AHEAD_POLY[1023-32* 30 -18])^(c[19]&AHEAD_POLY[1023-32* 30 -19])^(c[20]&AHEAD_POLY[1023-32* 30 -20])^(c[21]&AHEAD_POLY[1023-32* 30 -21])^(c[22]&AHEAD_POLY[1023-32* 30 -22])^(c[23]&AHEAD_POLY[1023-32* 30 -23])^(c[24]&AHEAD_POLY[1023-32* 30 -24])^(c[25]&AHEAD_POLY[1023-32* 30 -25])^(c[26]&AHEAD_POLY[1023-32* 30 -26])^(c[27]&AHEAD_POLY[1023-32* 30 -27])^(c[28]&AHEAD_POLY[1023-32* 30 -28])^(c[29]&AHEAD_POLY[1023-32* 30 -29])^(c[30]&AHEAD_POLY[1023-32* 30 -30])^(c[31]&AHEAD_POLY[1023-32* 30 -31]);
  //   newcrc[31]  = (c[0]&AHEAD_POLY[1023-32* 31 ])^(c[1]&AHEAD_POLY[1023-32* 31 -1])^(c[2]&AHEAD_POLY[1023-32* -2 ])^(c[3]&AHEAD_POLY[1023-32* 31 -3])^(c[4]&AHEAD_POLY[1023-32* 31 -4])^(c[5]&AHEAD_POLY[1023-32* 31 -5])^(c[6]&AHEAD_POLY[1023-32* 31 -6])^(c[7]&AHEAD_POLY[1023-32* 31 -7])^(c[8]&AHEAD_POLY[1023-32* 31 -8])^(c[9]&AHEAD_POLY[1023-32* 31 -9])^(c[10]&AHEAD_POLY[1023-32* 31 -10])^(c[11]&AHEAD_POLY[1023-32* 31 -11])^(c[12]&AHEAD_POLY[1023-32* 31 -12])^(c[13]&AHEAD_POLY[1023-32* 31 -13])^(c[14]&AHEAD_POLY[1023-32* 31 -14])^(c[15]&AHEAD_POLY[1023-32* 31 -15])^(c[16]&AHEAD_POLY[1023-32* 31 -16])^(c[17]&AHEAD_POLY[1023-32* 31 -17])^(c[18]&AHEAD_POLY[1023-32* 31 -18])^(c[19]&AHEAD_POLY[1023-32* 31 -19])^(c[20]&AHEAD_POLY[1023-32* 31 -20])^(c[21]&AHEAD_POLY[1023-32* 31 -21])^(c[22]&AHEAD_POLY[1023-32* 31 -22])^(c[23]&AHEAD_POLY[1023-32* 31 -23])^(c[24]&AHEAD_POLY[1023-32* 31 -24])^(c[25]&AHEAD_POLY[1023-32* 31 -25])^(c[26]&AHEAD_POLY[1023-32* 31 -26])^(c[27]&AHEAD_POLY[1023-32* 31 -27])^(c[28]&AHEAD_POLY[1023-32* 31 -28])^(c[29]&AHEAD_POLY[1023-32* 31 -29])^(c[30]&AHEAD_POLY[1023-32* 31 -30])^(c[31]&AHEAD_POLY[1023-32* 31 -31]);
  //   CRC32_ahead = newcrc;
  // end
  // endfunction


  //  function [31:0] CRC32_ahead;

  //   input [31:0] crc_i;
  //   // input [31:0] crc_o;
  //   //reg [31:0] d;
  //   reg [31:0] c;
  //   reg [31:0] newcrc;
  // begin
  //   c = crc_i;

  //   newcrc[0 ]  = (c[0]&ahead[1023-32* 0  ])^(c[1]&ahead[1023-32* 0  -1])^(c[2]&ahead[1023-32* -2 ])^(c[3]&ahead[1023-32* 0  -3])^(c[4]&ahead[1023-32* 0  -4])^(c[5]&ahead[1023-32* 0  -5])^(c[6]&ahead[1023-32* 0  -6])^(c[7]&ahead[1023-32* 0  -7])^(c[8]&ahead[1023-32* 0  -8])^(c[9]&ahead[1023-32* 0  -9])^(c[10]&ahead[1023-32* 0  -10])^(c[11]&ahead[1023-32* 0  -11])^(c[12]&ahead[1023-32* 0  -12])^(c[13]&ahead[1023-32* 0  -13])^(c[14]&ahead[1023-32* 0  -14])^(c[15]&ahead[1023-32* 0  -15])^(c[16]&ahead[1023-32* 0  -16])^(c[17]&ahead[1023-32* 0  -17])^(c[18]&ahead[1023-32* 0  -18])^(c[19]&ahead[1023-32* 0  -19])^(c[20]&ahead[1023-32* 0  -20])^(c[21]&ahead[1023-32* 0  -21])^(c[22]&ahead[1023-32* 0  -22])^(c[23]&ahead[1023-32* 0  -23])^(c[24]&ahead[1023-32* 0  -24])^(c[25]&ahead[1023-32* 0  -25])^(c[26]&ahead[1023-32* 0  -26])^(c[27]&ahead[1023-32* 0  -27])^(c[28]&ahead[1023-32* 0  -28])^(c[29]&ahead[1023-32* 0  -29])^(c[30]&ahead[1023-32* 0  -30])^(c[31]&ahead[1023-32* 0  -31]);
  //   newcrc[1 ]  = (c[0]&ahead[1023-32* 1  ])^(c[1]&ahead[1023-32* 1  -1])^(c[2]&ahead[1023-32* -2 ])^(c[3]&ahead[1023-32* 1  -3])^(c[4]&ahead[1023-32* 1  -4])^(c[5]&ahead[1023-32* 1  -5])^(c[6]&ahead[1023-32* 1  -6])^(c[7]&ahead[1023-32* 1  -7])^(c[8]&ahead[1023-32* 1  -8])^(c[9]&ahead[1023-32* 1  -9])^(c[10]&ahead[1023-32* 1  -10])^(c[11]&ahead[1023-32* 1  -11])^(c[12]&ahead[1023-32* 1  -12])^(c[13]&ahead[1023-32* 1  -13])^(c[14]&ahead[1023-32* 1  -14])^(c[15]&ahead[1023-32* 1  -15])^(c[16]&ahead[1023-32* 1  -16])^(c[17]&ahead[1023-32* 1  -17])^(c[18]&ahead[1023-32* 1  -18])^(c[19]&ahead[1023-32* 1  -19])^(c[20]&ahead[1023-32* 1  -20])^(c[21]&ahead[1023-32* 1  -21])^(c[22]&ahead[1023-32* 1  -22])^(c[23]&ahead[1023-32* 1  -23])^(c[24]&ahead[1023-32* 1  -24])^(c[25]&ahead[1023-32* 1  -25])^(c[26]&ahead[1023-32* 1  -26])^(c[27]&ahead[1023-32* 1  -27])^(c[28]&ahead[1023-32* 1  -28])^(c[29]&ahead[1023-32* 1  -29])^(c[30]&ahead[1023-32* 1  -30])^(c[31]&ahead[1023-32* 1  -31]);
  //   newcrc[2 ]  = (c[0]&ahead[1023-32* 2  ])^(c[1]&ahead[1023-32* 2  -1])^(c[2]&ahead[1023-32* -2 ])^(c[3]&ahead[1023-32* 2  -3])^(c[4]&ahead[1023-32* 2  -4])^(c[5]&ahead[1023-32* 2  -5])^(c[6]&ahead[1023-32* 2  -6])^(c[7]&ahead[1023-32* 2  -7])^(c[8]&ahead[1023-32* 2  -8])^(c[9]&ahead[1023-32* 2  -9])^(c[10]&ahead[1023-32* 2  -10])^(c[11]&ahead[1023-32* 2  -11])^(c[12]&ahead[1023-32* 2  -12])^(c[13]&ahead[1023-32* 2  -13])^(c[14]&ahead[1023-32* 2  -14])^(c[15]&ahead[1023-32* 2  -15])^(c[16]&ahead[1023-32* 2  -16])^(c[17]&ahead[1023-32* 2  -17])^(c[18]&ahead[1023-32* 2  -18])^(c[19]&ahead[1023-32* 2  -19])^(c[20]&ahead[1023-32* 2  -20])^(c[21]&ahead[1023-32* 2  -21])^(c[22]&ahead[1023-32* 2  -22])^(c[23]&ahead[1023-32* 2  -23])^(c[24]&ahead[1023-32* 2  -24])^(c[25]&ahead[1023-32* 2  -25])^(c[26]&ahead[1023-32* 2  -26])^(c[27]&ahead[1023-32* 2  -27])^(c[28]&ahead[1023-32* 2  -28])^(c[29]&ahead[1023-32* 2  -29])^(c[30]&ahead[1023-32* 2  -30])^(c[31]&ahead[1023-32* 2  -31]);
  //   newcrc[3 ]  = (c[0]&ahead[1023-32* 3  ])^(c[1]&ahead[1023-32* 3  -1])^(c[2]&ahead[1023-32* -2 ])^(c[3]&ahead[1023-32* 3  -3])^(c[4]&ahead[1023-32* 3  -4])^(c[5]&ahead[1023-32* 3  -5])^(c[6]&ahead[1023-32* 3  -6])^(c[7]&ahead[1023-32* 3  -7])^(c[8]&ahead[1023-32* 3  -8])^(c[9]&ahead[1023-32* 3  -9])^(c[10]&ahead[1023-32* 3  -10])^(c[11]&ahead[1023-32* 3  -11])^(c[12]&ahead[1023-32* 3  -12])^(c[13]&ahead[1023-32* 3  -13])^(c[14]&ahead[1023-32* 3  -14])^(c[15]&ahead[1023-32* 3  -15])^(c[16]&ahead[1023-32* 3  -16])^(c[17]&ahead[1023-32* 3  -17])^(c[18]&ahead[1023-32* 3  -18])^(c[19]&ahead[1023-32* 3  -19])^(c[20]&ahead[1023-32* 3  -20])^(c[21]&ahead[1023-32* 3  -21])^(c[22]&ahead[1023-32* 3  -22])^(c[23]&ahead[1023-32* 3  -23])^(c[24]&ahead[1023-32* 3  -24])^(c[25]&ahead[1023-32* 3  -25])^(c[26]&ahead[1023-32* 3  -26])^(c[27]&ahead[1023-32* 3  -27])^(c[28]&ahead[1023-32* 3  -28])^(c[29]&ahead[1023-32* 3  -29])^(c[30]&ahead[1023-32* 3  -30])^(c[31]&ahead[1023-32* 3  -31]);
  //   newcrc[4 ]  = (c[0]&ahead[1023-32* 4  ])^(c[1]&ahead[1023-32* 4  -1])^(c[2]&ahead[1023-32* -2 ])^(c[3]&ahead[1023-32* 4  -3])^(c[4]&ahead[1023-32* 4  -4])^(c[5]&ahead[1023-32* 4  -5])^(c[6]&ahead[1023-32* 4  -6])^(c[7]&ahead[1023-32* 4  -7])^(c[8]&ahead[1023-32* 4  -8])^(c[9]&ahead[1023-32* 4  -9])^(c[10]&ahead[1023-32* 4  -10])^(c[11]&ahead[1023-32* 4  -11])^(c[12]&ahead[1023-32* 4  -12])^(c[13]&ahead[1023-32* 4  -13])^(c[14]&ahead[1023-32* 4  -14])^(c[15]&ahead[1023-32* 4  -15])^(c[16]&ahead[1023-32* 4  -16])^(c[17]&ahead[1023-32* 4  -17])^(c[18]&ahead[1023-32* 4  -18])^(c[19]&ahead[1023-32* 4  -19])^(c[20]&ahead[1023-32* 4  -20])^(c[21]&ahead[1023-32* 4  -21])^(c[22]&ahead[1023-32* 4  -22])^(c[23]&ahead[1023-32* 4  -23])^(c[24]&ahead[1023-32* 4  -24])^(c[25]&ahead[1023-32* 4  -25])^(c[26]&ahead[1023-32* 4  -26])^(c[27]&ahead[1023-32* 4  -27])^(c[28]&ahead[1023-32* 4  -28])^(c[29]&ahead[1023-32* 4  -29])^(c[30]&ahead[1023-32* 4  -30])^(c[31]&ahead[1023-32* 4  -31]);
  //   newcrc[5 ]  = (c[0]&ahead[1023-32* 5  ])^(c[1]&ahead[1023-32* 5  -1])^(c[2]&ahead[1023-32* -2 ])^(c[3]&ahead[1023-32* 5  -3])^(c[4]&ahead[1023-32* 5  -4])^(c[5]&ahead[1023-32* 5  -5])^(c[6]&ahead[1023-32* 5  -6])^(c[7]&ahead[1023-32* 5  -7])^(c[8]&ahead[1023-32* 5  -8])^(c[9]&ahead[1023-32* 5  -9])^(c[10]&ahead[1023-32* 5  -10])^(c[11]&ahead[1023-32* 5  -11])^(c[12]&ahead[1023-32* 5  -12])^(c[13]&ahead[1023-32* 5  -13])^(c[14]&ahead[1023-32* 5  -14])^(c[15]&ahead[1023-32* 5  -15])^(c[16]&ahead[1023-32* 5  -16])^(c[17]&ahead[1023-32* 5  -17])^(c[18]&ahead[1023-32* 5  -18])^(c[19]&ahead[1023-32* 5  -19])^(c[20]&ahead[1023-32* 5  -20])^(c[21]&ahead[1023-32* 5  -21])^(c[22]&ahead[1023-32* 5  -22])^(c[23]&ahead[1023-32* 5  -23])^(c[24]&ahead[1023-32* 5  -24])^(c[25]&ahead[1023-32* 5  -25])^(c[26]&ahead[1023-32* 5  -26])^(c[27]&ahead[1023-32* 5  -27])^(c[28]&ahead[1023-32* 5  -28])^(c[29]&ahead[1023-32* 5  -29])^(c[30]&ahead[1023-32* 5  -30])^(c[31]&ahead[1023-32* 5  -31]);
  //   newcrc[6 ]  = (c[0]&ahead[1023-32* 6  ])^(c[1]&ahead[1023-32* 6  -1])^(c[2]&ahead[1023-32* -2 ])^(c[3]&ahead[1023-32* 6  -3])^(c[4]&ahead[1023-32* 6  -4])^(c[5]&ahead[1023-32* 6  -5])^(c[6]&ahead[1023-32* 6  -6])^(c[7]&ahead[1023-32* 6  -7])^(c[8]&ahead[1023-32* 6  -8])^(c[9]&ahead[1023-32* 6  -9])^(c[10]&ahead[1023-32* 6  -10])^(c[11]&ahead[1023-32* 6  -11])^(c[12]&ahead[1023-32* 6  -12])^(c[13]&ahead[1023-32* 6  -13])^(c[14]&ahead[1023-32* 6  -14])^(c[15]&ahead[1023-32* 6  -15])^(c[16]&ahead[1023-32* 6  -16])^(c[17]&ahead[1023-32* 6  -17])^(c[18]&ahead[1023-32* 6  -18])^(c[19]&ahead[1023-32* 6  -19])^(c[20]&ahead[1023-32* 6  -20])^(c[21]&ahead[1023-32* 6  -21])^(c[22]&ahead[1023-32* 6  -22])^(c[23]&ahead[1023-32* 6  -23])^(c[24]&ahead[1023-32* 6  -24])^(c[25]&ahead[1023-32* 6  -25])^(c[26]&ahead[1023-32* 6  -26])^(c[27]&ahead[1023-32* 6  -27])^(c[28]&ahead[1023-32* 6  -28])^(c[29]&ahead[1023-32* 6  -29])^(c[30]&ahead[1023-32* 6  -30])^(c[31]&ahead[1023-32* 6  -31]);
  //   newcrc[7 ]  = (c[0]&ahead[1023-32* 7  ])^(c[1]&ahead[1023-32* 7  -1])^(c[2]&ahead[1023-32* -2 ])^(c[3]&ahead[1023-32* 7  -3])^(c[4]&ahead[1023-32* 7  -4])^(c[5]&ahead[1023-32* 7  -5])^(c[6]&ahead[1023-32* 7  -6])^(c[7]&ahead[1023-32* 7  -7])^(c[8]&ahead[1023-32* 7  -8])^(c[9]&ahead[1023-32* 7  -9])^(c[10]&ahead[1023-32* 7  -10])^(c[11]&ahead[1023-32* 7  -11])^(c[12]&ahead[1023-32* 7  -12])^(c[13]&ahead[1023-32* 7  -13])^(c[14]&ahead[1023-32* 7  -14])^(c[15]&ahead[1023-32* 7  -15])^(c[16]&ahead[1023-32* 7  -16])^(c[17]&ahead[1023-32* 7  -17])^(c[18]&ahead[1023-32* 7  -18])^(c[19]&ahead[1023-32* 7  -19])^(c[20]&ahead[1023-32* 7  -20])^(c[21]&ahead[1023-32* 7  -21])^(c[22]&ahead[1023-32* 7  -22])^(c[23]&ahead[1023-32* 7  -23])^(c[24]&ahead[1023-32* 7  -24])^(c[25]&ahead[1023-32* 7  -25])^(c[26]&ahead[1023-32* 7  -26])^(c[27]&ahead[1023-32* 7  -27])^(c[28]&ahead[1023-32* 7  -28])^(c[29]&ahead[1023-32* 7  -29])^(c[30]&ahead[1023-32* 7  -30])^(c[31]&ahead[1023-32* 7  -31]);
  //   newcrc[8 ]  = (c[0]&ahead[1023-32* 8  ])^(c[1]&ahead[1023-32* 8  -1])^(c[2]&ahead[1023-32* -2 ])^(c[3]&ahead[1023-32* 8  -3])^(c[4]&ahead[1023-32* 8  -4])^(c[5]&ahead[1023-32* 8  -5])^(c[6]&ahead[1023-32* 8  -6])^(c[7]&ahead[1023-32* 8  -7])^(c[8]&ahead[1023-32* 8  -8])^(c[9]&ahead[1023-32* 8  -9])^(c[10]&ahead[1023-32* 8  -10])^(c[11]&ahead[1023-32* 8  -11])^(c[12]&ahead[1023-32* 8  -12])^(c[13]&ahead[1023-32* 8  -13])^(c[14]&ahead[1023-32* 8  -14])^(c[15]&ahead[1023-32* 8  -15])^(c[16]&ahead[1023-32* 8  -16])^(c[17]&ahead[1023-32* 8  -17])^(c[18]&ahead[1023-32* 8  -18])^(c[19]&ahead[1023-32* 8  -19])^(c[20]&ahead[1023-32* 8  -20])^(c[21]&ahead[1023-32* 8  -21])^(c[22]&ahead[1023-32* 8  -22])^(c[23]&ahead[1023-32* 8  -23])^(c[24]&ahead[1023-32* 8  -24])^(c[25]&ahead[1023-32* 8  -25])^(c[26]&ahead[1023-32* 8  -26])^(c[27]&ahead[1023-32* 8  -27])^(c[28]&ahead[1023-32* 8  -28])^(c[29]&ahead[1023-32* 8  -29])^(c[30]&ahead[1023-32* 8  -30])^(c[31]&ahead[1023-32* 8  -31]);
  //   newcrc[9 ]  = (c[0]&ahead[1023-32* 9  ])^(c[1]&ahead[1023-32* 9  -1])^(c[2]&ahead[1023-32* -2 ])^(c[3]&ahead[1023-32* 9  -3])^(c[4]&ahead[1023-32* 9  -4])^(c[5]&ahead[1023-32* 9  -5])^(c[6]&ahead[1023-32* 9  -6])^(c[7]&ahead[1023-32* 9  -7])^(c[8]&ahead[1023-32* 9  -8])^(c[9]&ahead[1023-32* 9  -9])^(c[10]&ahead[1023-32* 9  -10])^(c[11]&ahead[1023-32* 9  -11])^(c[12]&ahead[1023-32* 9  -12])^(c[13]&ahead[1023-32* 9  -13])^(c[14]&ahead[1023-32* 9  -14])^(c[15]&ahead[1023-32* 9  -15])^(c[16]&ahead[1023-32* 9  -16])^(c[17]&ahead[1023-32* 9  -17])^(c[18]&ahead[1023-32* 9  -18])^(c[19]&ahead[1023-32* 9  -19])^(c[20]&ahead[1023-32* 9  -20])^(c[21]&ahead[1023-32* 9  -21])^(c[22]&ahead[1023-32* 9  -22])^(c[23]&ahead[1023-32* 9  -23])^(c[24]&ahead[1023-32* 9  -24])^(c[25]&ahead[1023-32* 9  -25])^(c[26]&ahead[1023-32* 9  -26])^(c[27]&ahead[1023-32* 9  -27])^(c[28]&ahead[1023-32* 9  -28])^(c[29]&ahead[1023-32* 9  -29])^(c[30]&ahead[1023-32* 9  -30])^(c[31]&ahead[1023-32* 9  -31]);
  //   newcrc[10]  = (c[0]&ahead[1023-32* 10 ])^(c[1]&ahead[1023-32* 10 -1])^(c[2]&ahead[1023-32* -2 ])^(c[3]&ahead[1023-32* 10 -3])^(c[4]&ahead[1023-32* 10 -4])^(c[5]&ahead[1023-32* 10 -5])^(c[6]&ahead[1023-32* 10 -6])^(c[7]&ahead[1023-32* 10 -7])^(c[8]&ahead[1023-32* 10 -8])^(c[9]&ahead[1023-32* 10 -9])^(c[10]&ahead[1023-32* 10 -10])^(c[11]&ahead[1023-32* 10 -11])^(c[12]&ahead[1023-32* 10 -12])^(c[13]&ahead[1023-32* 10 -13])^(c[14]&ahead[1023-32* 10 -14])^(c[15]&ahead[1023-32* 10 -15])^(c[16]&ahead[1023-32* 10 -16])^(c[17]&ahead[1023-32* 10 -17])^(c[18]&ahead[1023-32* 10 -18])^(c[19]&ahead[1023-32* 10 -19])^(c[20]&ahead[1023-32* 10 -20])^(c[21]&ahead[1023-32* 10 -21])^(c[22]&ahead[1023-32* 10 -22])^(c[23]&ahead[1023-32* 10 -23])^(c[24]&ahead[1023-32* 10 -24])^(c[25]&ahead[1023-32* 10 -25])^(c[26]&ahead[1023-32* 10 -26])^(c[27]&ahead[1023-32* 10 -27])^(c[28]&ahead[1023-32* 10 -28])^(c[29]&ahead[1023-32* 10 -29])^(c[30]&ahead[1023-32* 10 -30])^(c[31]&ahead[1023-32* 10 -31]);
  //   newcrc[11]  = (c[0]&ahead[1023-32* 11 ])^(c[1]&ahead[1023-32* 11 -1])^(c[2]&ahead[1023-32* -2 ])^(c[3]&ahead[1023-32* 11 -3])^(c[4]&ahead[1023-32* 11 -4])^(c[5]&ahead[1023-32* 11 -5])^(c[6]&ahead[1023-32* 11 -6])^(c[7]&ahead[1023-32* 11 -7])^(c[8]&ahead[1023-32* 11 -8])^(c[9]&ahead[1023-32* 11 -9])^(c[10]&ahead[1023-32* 11 -10])^(c[11]&ahead[1023-32* 11 -11])^(c[12]&ahead[1023-32* 11 -12])^(c[13]&ahead[1023-32* 11 -13])^(c[14]&ahead[1023-32* 11 -14])^(c[15]&ahead[1023-32* 11 -15])^(c[16]&ahead[1023-32* 11 -16])^(c[17]&ahead[1023-32* 11 -17])^(c[18]&ahead[1023-32* 11 -18])^(c[19]&ahead[1023-32* 11 -19])^(c[20]&ahead[1023-32* 11 -20])^(c[21]&ahead[1023-32* 11 -21])^(c[22]&ahead[1023-32* 11 -22])^(c[23]&ahead[1023-32* 11 -23])^(c[24]&ahead[1023-32* 11 -24])^(c[25]&ahead[1023-32* 11 -25])^(c[26]&ahead[1023-32* 11 -26])^(c[27]&ahead[1023-32* 11 -27])^(c[28]&ahead[1023-32* 11 -28])^(c[29]&ahead[1023-32* 11 -29])^(c[30]&ahead[1023-32* 11 -30])^(c[31]&ahead[1023-32* 11 -31]);
  //   newcrc[12]  = (c[0]&ahead[1023-32* 12 ])^(c[1]&ahead[1023-32* 12 -1])^(c[2]&ahead[1023-32* -2 ])^(c[3]&ahead[1023-32* 12 -3])^(c[4]&ahead[1023-32* 12 -4])^(c[5]&ahead[1023-32* 12 -5])^(c[6]&ahead[1023-32* 12 -6])^(c[7]&ahead[1023-32* 12 -7])^(c[8]&ahead[1023-32* 12 -8])^(c[9]&ahead[1023-32* 12 -9])^(c[10]&ahead[1023-32* 12 -10])^(c[11]&ahead[1023-32* 12 -11])^(c[12]&ahead[1023-32* 12 -12])^(c[13]&ahead[1023-32* 12 -13])^(c[14]&ahead[1023-32* 12 -14])^(c[15]&ahead[1023-32* 12 -15])^(c[16]&ahead[1023-32* 12 -16])^(c[17]&ahead[1023-32* 12 -17])^(c[18]&ahead[1023-32* 12 -18])^(c[19]&ahead[1023-32* 12 -19])^(c[20]&ahead[1023-32* 12 -20])^(c[21]&ahead[1023-32* 12 -21])^(c[22]&ahead[1023-32* 12 -22])^(c[23]&ahead[1023-32* 12 -23])^(c[24]&ahead[1023-32* 12 -24])^(c[25]&ahead[1023-32* 12 -25])^(c[26]&ahead[1023-32* 12 -26])^(c[27]&ahead[1023-32* 12 -27])^(c[28]&ahead[1023-32* 12 -28])^(c[29]&ahead[1023-32* 12 -29])^(c[30]&ahead[1023-32* 12 -30])^(c[31]&ahead[1023-32* 12 -31]);
  //   newcrc[13]  = (c[0]&ahead[1023-32* 13 ])^(c[1]&ahead[1023-32* 13 -1])^(c[2]&ahead[1023-32* -2 ])^(c[3]&ahead[1023-32* 13 -3])^(c[4]&ahead[1023-32* 13 -4])^(c[5]&ahead[1023-32* 13 -5])^(c[6]&ahead[1023-32* 13 -6])^(c[7]&ahead[1023-32* 13 -7])^(c[8]&ahead[1023-32* 13 -8])^(c[9]&ahead[1023-32* 13 -9])^(c[10]&ahead[1023-32* 13 -10])^(c[11]&ahead[1023-32* 13 -11])^(c[12]&ahead[1023-32* 13 -12])^(c[13]&ahead[1023-32* 13 -13])^(c[14]&ahead[1023-32* 13 -14])^(c[15]&ahead[1023-32* 13 -15])^(c[16]&ahead[1023-32* 13 -16])^(c[17]&ahead[1023-32* 13 -17])^(c[18]&ahead[1023-32* 13 -18])^(c[19]&ahead[1023-32* 13 -19])^(c[20]&ahead[1023-32* 13 -20])^(c[21]&ahead[1023-32* 13 -21])^(c[22]&ahead[1023-32* 13 -22])^(c[23]&ahead[1023-32* 13 -23])^(c[24]&ahead[1023-32* 13 -24])^(c[25]&ahead[1023-32* 13 -25])^(c[26]&ahead[1023-32* 13 -26])^(c[27]&ahead[1023-32* 13 -27])^(c[28]&ahead[1023-32* 13 -28])^(c[29]&ahead[1023-32* 13 -29])^(c[30]&ahead[1023-32* 13 -30])^(c[31]&ahead[1023-32* 13 -31]);
  //   newcrc[14]  = (c[0]&ahead[1023-32* 14 ])^(c[1]&ahead[1023-32* 14 -1])^(c[2]&ahead[1023-32* -2 ])^(c[3]&ahead[1023-32* 14 -3])^(c[4]&ahead[1023-32* 14 -4])^(c[5]&ahead[1023-32* 14 -5])^(c[6]&ahead[1023-32* 14 -6])^(c[7]&ahead[1023-32* 14 -7])^(c[8]&ahead[1023-32* 14 -8])^(c[9]&ahead[1023-32* 14 -9])^(c[10]&ahead[1023-32* 14 -10])^(c[11]&ahead[1023-32* 14 -11])^(c[12]&ahead[1023-32* 14 -12])^(c[13]&ahead[1023-32* 14 -13])^(c[14]&ahead[1023-32* 14 -14])^(c[15]&ahead[1023-32* 14 -15])^(c[16]&ahead[1023-32* 14 -16])^(c[17]&ahead[1023-32* 14 -17])^(c[18]&ahead[1023-32* 14 -18])^(c[19]&ahead[1023-32* 14 -19])^(c[20]&ahead[1023-32* 14 -20])^(c[21]&ahead[1023-32* 14 -21])^(c[22]&ahead[1023-32* 14 -22])^(c[23]&ahead[1023-32* 14 -23])^(c[24]&ahead[1023-32* 14 -24])^(c[25]&ahead[1023-32* 14 -25])^(c[26]&ahead[1023-32* 14 -26])^(c[27]&ahead[1023-32* 14 -27])^(c[28]&ahead[1023-32* 14 -28])^(c[29]&ahead[1023-32* 14 -29])^(c[30]&ahead[1023-32* 14 -30])^(c[31]&ahead[1023-32* 14 -31]);
  //   newcrc[15]  = (c[0]&ahead[1023-32* 15 ])^(c[1]&ahead[1023-32* 15 -1])^(c[2]&ahead[1023-32* -2 ])^(c[3]&ahead[1023-32* 15 -3])^(c[4]&ahead[1023-32* 15 -4])^(c[5]&ahead[1023-32* 15 -5])^(c[6]&ahead[1023-32* 15 -6])^(c[7]&ahead[1023-32* 15 -7])^(c[8]&ahead[1023-32* 15 -8])^(c[9]&ahead[1023-32* 15 -9])^(c[10]&ahead[1023-32* 15 -10])^(c[11]&ahead[1023-32* 15 -11])^(c[12]&ahead[1023-32* 15 -12])^(c[13]&ahead[1023-32* 15 -13])^(c[14]&ahead[1023-32* 15 -14])^(c[15]&ahead[1023-32* 15 -15])^(c[16]&ahead[1023-32* 15 -16])^(c[17]&ahead[1023-32* 15 -17])^(c[18]&ahead[1023-32* 15 -18])^(c[19]&ahead[1023-32* 15 -19])^(c[20]&ahead[1023-32* 15 -20])^(c[21]&ahead[1023-32* 15 -21])^(c[22]&ahead[1023-32* 15 -22])^(c[23]&ahead[1023-32* 15 -23])^(c[24]&ahead[1023-32* 15 -24])^(c[25]&ahead[1023-32* 15 -25])^(c[26]&ahead[1023-32* 15 -26])^(c[27]&ahead[1023-32* 15 -27])^(c[28]&ahead[1023-32* 15 -28])^(c[29]&ahead[1023-32* 15 -29])^(c[30]&ahead[1023-32* 15 -30])^(c[31]&ahead[1023-32* 15 -31]);
  //   newcrc[16]  = (c[0]&ahead[1023-32* 16 ])^(c[1]&ahead[1023-32* 16 -1])^(c[2]&ahead[1023-32* -2 ])^(c[3]&ahead[1023-32* 16 -3])^(c[4]&ahead[1023-32* 16 -4])^(c[5]&ahead[1023-32* 16 -5])^(c[6]&ahead[1023-32* 16 -6])^(c[7]&ahead[1023-32* 16 -7])^(c[8]&ahead[1023-32* 16 -8])^(c[9]&ahead[1023-32* 16 -9])^(c[10]&ahead[1023-32* 16 -10])^(c[11]&ahead[1023-32* 16 -11])^(c[12]&ahead[1023-32* 16 -12])^(c[13]&ahead[1023-32* 16 -13])^(c[14]&ahead[1023-32* 16 -14])^(c[15]&ahead[1023-32* 16 -15])^(c[16]&ahead[1023-32* 16 -16])^(c[17]&ahead[1023-32* 16 -17])^(c[18]&ahead[1023-32* 16 -18])^(c[19]&ahead[1023-32* 16 -19])^(c[20]&ahead[1023-32* 16 -20])^(c[21]&ahead[1023-32* 16 -21])^(c[22]&ahead[1023-32* 16 -22])^(c[23]&ahead[1023-32* 16 -23])^(c[24]&ahead[1023-32* 16 -24])^(c[25]&ahead[1023-32* 16 -25])^(c[26]&ahead[1023-32* 16 -26])^(c[27]&ahead[1023-32* 16 -27])^(c[28]&ahead[1023-32* 16 -28])^(c[29]&ahead[1023-32* 16 -29])^(c[30]&ahead[1023-32* 16 -30])^(c[31]&ahead[1023-32* 16 -31]);
  //   newcrc[17]  = (c[0]&ahead[1023-32* 17 ])^(c[1]&ahead[1023-32* 17 -1])^(c[2]&ahead[1023-32* -2 ])^(c[3]&ahead[1023-32* 17 -3])^(c[4]&ahead[1023-32* 17 -4])^(c[5]&ahead[1023-32* 17 -5])^(c[6]&ahead[1023-32* 17 -6])^(c[7]&ahead[1023-32* 17 -7])^(c[8]&ahead[1023-32* 17 -8])^(c[9]&ahead[1023-32* 17 -9])^(c[10]&ahead[1023-32* 17 -10])^(c[11]&ahead[1023-32* 17 -11])^(c[12]&ahead[1023-32* 17 -12])^(c[13]&ahead[1023-32* 17 -13])^(c[14]&ahead[1023-32* 17 -14])^(c[15]&ahead[1023-32* 17 -15])^(c[16]&ahead[1023-32* 17 -16])^(c[17]&ahead[1023-32* 17 -17])^(c[18]&ahead[1023-32* 17 -18])^(c[19]&ahead[1023-32* 17 -19])^(c[20]&ahead[1023-32* 17 -20])^(c[21]&ahead[1023-32* 17 -21])^(c[22]&ahead[1023-32* 17 -22])^(c[23]&ahead[1023-32* 17 -23])^(c[24]&ahead[1023-32* 17 -24])^(c[25]&ahead[1023-32* 17 -25])^(c[26]&ahead[1023-32* 17 -26])^(c[27]&ahead[1023-32* 17 -27])^(c[28]&ahead[1023-32* 17 -28])^(c[29]&ahead[1023-32* 17 -29])^(c[30]&ahead[1023-32* 17 -30])^(c[31]&ahead[1023-32* 17 -31]);
  //   newcrc[18]  = (c[0]&ahead[1023-32* 18 ])^(c[1]&ahead[1023-32* 18 -1])^(c[2]&ahead[1023-32* -2 ])^(c[3]&ahead[1023-32* 18 -3])^(c[4]&ahead[1023-32* 18 -4])^(c[5]&ahead[1023-32* 18 -5])^(c[6]&ahead[1023-32* 18 -6])^(c[7]&ahead[1023-32* 18 -7])^(c[8]&ahead[1023-32* 18 -8])^(c[9]&ahead[1023-32* 18 -9])^(c[10]&ahead[1023-32* 18 -10])^(c[11]&ahead[1023-32* 18 -11])^(c[12]&ahead[1023-32* 18 -12])^(c[13]&ahead[1023-32* 18 -13])^(c[14]&ahead[1023-32* 18 -14])^(c[15]&ahead[1023-32* 18 -15])^(c[16]&ahead[1023-32* 18 -16])^(c[17]&ahead[1023-32* 18 -17])^(c[18]&ahead[1023-32* 18 -18])^(c[19]&ahead[1023-32* 18 -19])^(c[20]&ahead[1023-32* 18 -20])^(c[21]&ahead[1023-32* 18 -21])^(c[22]&ahead[1023-32* 18 -22])^(c[23]&ahead[1023-32* 18 -23])^(c[24]&ahead[1023-32* 18 -24])^(c[25]&ahead[1023-32* 18 -25])^(c[26]&ahead[1023-32* 18 -26])^(c[27]&ahead[1023-32* 18 -27])^(c[28]&ahead[1023-32* 18 -28])^(c[29]&ahead[1023-32* 18 -29])^(c[30]&ahead[1023-32* 18 -30])^(c[31]&ahead[1023-32* 18 -31]);
  //   newcrc[19]  = (c[0]&ahead[1023-32* 19 ])^(c[1]&ahead[1023-32* 19 -1])^(c[2]&ahead[1023-32* -2 ])^(c[3]&ahead[1023-32* 19 -3])^(c[4]&ahead[1023-32* 19 -4])^(c[5]&ahead[1023-32* 19 -5])^(c[6]&ahead[1023-32* 19 -6])^(c[7]&ahead[1023-32* 19 -7])^(c[8]&ahead[1023-32* 19 -8])^(c[9]&ahead[1023-32* 19 -9])^(c[10]&ahead[1023-32* 19 -10])^(c[11]&ahead[1023-32* 19 -11])^(c[12]&ahead[1023-32* 19 -12])^(c[13]&ahead[1023-32* 19 -13])^(c[14]&ahead[1023-32* 19 -14])^(c[15]&ahead[1023-32* 19 -15])^(c[16]&ahead[1023-32* 19 -16])^(c[17]&ahead[1023-32* 19 -17])^(c[18]&ahead[1023-32* 19 -18])^(c[19]&ahead[1023-32* 19 -19])^(c[20]&ahead[1023-32* 19 -20])^(c[21]&ahead[1023-32* 19 -21])^(c[22]&ahead[1023-32* 19 -22])^(c[23]&ahead[1023-32* 19 -23])^(c[24]&ahead[1023-32* 19 -24])^(c[25]&ahead[1023-32* 19 -25])^(c[26]&ahead[1023-32* 19 -26])^(c[27]&ahead[1023-32* 19 -27])^(c[28]&ahead[1023-32* 19 -28])^(c[29]&ahead[1023-32* 19 -29])^(c[30]&ahead[1023-32* 19 -30])^(c[31]&ahead[1023-32* 19 -31]);
  //   newcrc[20]  = (c[0]&ahead[1023-32* 20 ])^(c[1]&ahead[1023-32* 20 -1])^(c[2]&ahead[1023-32* -2 ])^(c[3]&ahead[1023-32* 20 -3])^(c[4]&ahead[1023-32* 20 -4])^(c[5]&ahead[1023-32* 20 -5])^(c[6]&ahead[1023-32* 20 -6])^(c[7]&ahead[1023-32* 20 -7])^(c[8]&ahead[1023-32* 20 -8])^(c[9]&ahead[1023-32* 20 -9])^(c[10]&ahead[1023-32* 20 -10])^(c[11]&ahead[1023-32* 20 -11])^(c[12]&ahead[1023-32* 20 -12])^(c[13]&ahead[1023-32* 20 -13])^(c[14]&ahead[1023-32* 20 -14])^(c[15]&ahead[1023-32* 20 -15])^(c[16]&ahead[1023-32* 20 -16])^(c[17]&ahead[1023-32* 20 -17])^(c[18]&ahead[1023-32* 20 -18])^(c[19]&ahead[1023-32* 20 -19])^(c[20]&ahead[1023-32* 20 -20])^(c[21]&ahead[1023-32* 20 -21])^(c[22]&ahead[1023-32* 20 -22])^(c[23]&ahead[1023-32* 20 -23])^(c[24]&ahead[1023-32* 20 -24])^(c[25]&ahead[1023-32* 20 -25])^(c[26]&ahead[1023-32* 20 -26])^(c[27]&ahead[1023-32* 20 -27])^(c[28]&ahead[1023-32* 20 -28])^(c[29]&ahead[1023-32* 20 -29])^(c[30]&ahead[1023-32* 20 -30])^(c[31]&ahead[1023-32* 20 -31]);
  //   newcrc[21]  = (c[0]&ahead[1023-32* 21 ])^(c[1]&ahead[1023-32* 21 -1])^(c[2]&ahead[1023-32* -2 ])^(c[3]&ahead[1023-32* 21 -3])^(c[4]&ahead[1023-32* 21 -4])^(c[5]&ahead[1023-32* 21 -5])^(c[6]&ahead[1023-32* 21 -6])^(c[7]&ahead[1023-32* 21 -7])^(c[8]&ahead[1023-32* 21 -8])^(c[9]&ahead[1023-32* 21 -9])^(c[10]&ahead[1023-32* 21 -10])^(c[11]&ahead[1023-32* 21 -11])^(c[12]&ahead[1023-32* 21 -12])^(c[13]&ahead[1023-32* 21 -13])^(c[14]&ahead[1023-32* 21 -14])^(c[15]&ahead[1023-32* 21 -15])^(c[16]&ahead[1023-32* 21 -16])^(c[17]&ahead[1023-32* 21 -17])^(c[18]&ahead[1023-32* 21 -18])^(c[19]&ahead[1023-32* 21 -19])^(c[20]&ahead[1023-32* 21 -20])^(c[21]&ahead[1023-32* 21 -21])^(c[22]&ahead[1023-32* 21 -22])^(c[23]&ahead[1023-32* 21 -23])^(c[24]&ahead[1023-32* 21 -24])^(c[25]&ahead[1023-32* 21 -25])^(c[26]&ahead[1023-32* 21 -26])^(c[27]&ahead[1023-32* 21 -27])^(c[28]&ahead[1023-32* 21 -28])^(c[29]&ahead[1023-32* 21 -29])^(c[30]&ahead[1023-32* 21 -30])^(c[31]&ahead[1023-32* 21 -31]);
  //   newcrc[22]  = (c[0]&ahead[1023-32* 22 ])^(c[1]&ahead[1023-32* 22 -1])^(c[2]&ahead[1023-32* -2 ])^(c[3]&ahead[1023-32* 22 -3])^(c[4]&ahead[1023-32* 22 -4])^(c[5]&ahead[1023-32* 22 -5])^(c[6]&ahead[1023-32* 22 -6])^(c[7]&ahead[1023-32* 22 -7])^(c[8]&ahead[1023-32* 22 -8])^(c[9]&ahead[1023-32* 22 -9])^(c[10]&ahead[1023-32* 22 -10])^(c[11]&ahead[1023-32* 22 -11])^(c[12]&ahead[1023-32* 22 -12])^(c[13]&ahead[1023-32* 22 -13])^(c[14]&ahead[1023-32* 22 -14])^(c[15]&ahead[1023-32* 22 -15])^(c[16]&ahead[1023-32* 22 -16])^(c[17]&ahead[1023-32* 22 -17])^(c[18]&ahead[1023-32* 22 -18])^(c[19]&ahead[1023-32* 22 -19])^(c[20]&ahead[1023-32* 22 -20])^(c[21]&ahead[1023-32* 22 -21])^(c[22]&ahead[1023-32* 22 -22])^(c[23]&ahead[1023-32* 22 -23])^(c[24]&ahead[1023-32* 22 -24])^(c[25]&ahead[1023-32* 22 -25])^(c[26]&ahead[1023-32* 22 -26])^(c[27]&ahead[1023-32* 22 -27])^(c[28]&ahead[1023-32* 22 -28])^(c[29]&ahead[1023-32* 22 -29])^(c[30]&ahead[1023-32* 22 -30])^(c[31]&ahead[1023-32* 22 -31]);
  //   newcrc[23]  = (c[0]&ahead[1023-32* 23 ])^(c[1]&ahead[1023-32* 23 -1])^(c[2]&ahead[1023-32* -2 ])^(c[3]&ahead[1023-32* 23 -3])^(c[4]&ahead[1023-32* 23 -4])^(c[5]&ahead[1023-32* 23 -5])^(c[6]&ahead[1023-32* 23 -6])^(c[7]&ahead[1023-32* 23 -7])^(c[8]&ahead[1023-32* 23 -8])^(c[9]&ahead[1023-32* 23 -9])^(c[10]&ahead[1023-32* 23 -10])^(c[11]&ahead[1023-32* 23 -11])^(c[12]&ahead[1023-32* 23 -12])^(c[13]&ahead[1023-32* 23 -13])^(c[14]&ahead[1023-32* 23 -14])^(c[15]&ahead[1023-32* 23 -15])^(c[16]&ahead[1023-32* 23 -16])^(c[17]&ahead[1023-32* 23 -17])^(c[18]&ahead[1023-32* 23 -18])^(c[19]&ahead[1023-32* 23 -19])^(c[20]&ahead[1023-32* 23 -20])^(c[21]&ahead[1023-32* 23 -21])^(c[22]&ahead[1023-32* 23 -22])^(c[23]&ahead[1023-32* 23 -23])^(c[24]&ahead[1023-32* 23 -24])^(c[25]&ahead[1023-32* 23 -25])^(c[26]&ahead[1023-32* 23 -26])^(c[27]&ahead[1023-32* 23 -27])^(c[28]&ahead[1023-32* 23 -28])^(c[29]&ahead[1023-32* 23 -29])^(c[30]&ahead[1023-32* 23 -30])^(c[31]&ahead[1023-32* 23 -31]);
  //   newcrc[24]  = (c[0]&ahead[1023-32* 24 ])^(c[1]&ahead[1023-32* 24 -1])^(c[2]&ahead[1023-32* -2 ])^(c[3]&ahead[1023-32* 24 -3])^(c[4]&ahead[1023-32* 24 -4])^(c[5]&ahead[1023-32* 24 -5])^(c[6]&ahead[1023-32* 24 -6])^(c[7]&ahead[1023-32* 24 -7])^(c[8]&ahead[1023-32* 24 -8])^(c[9]&ahead[1023-32* 24 -9])^(c[10]&ahead[1023-32* 24 -10])^(c[11]&ahead[1023-32* 24 -11])^(c[12]&ahead[1023-32* 24 -12])^(c[13]&ahead[1023-32* 24 -13])^(c[14]&ahead[1023-32* 24 -14])^(c[15]&ahead[1023-32* 24 -15])^(c[16]&ahead[1023-32* 24 -16])^(c[17]&ahead[1023-32* 24 -17])^(c[18]&ahead[1023-32* 24 -18])^(c[19]&ahead[1023-32* 24 -19])^(c[20]&ahead[1023-32* 24 -20])^(c[21]&ahead[1023-32* 24 -21])^(c[22]&ahead[1023-32* 24 -22])^(c[23]&ahead[1023-32* 24 -23])^(c[24]&ahead[1023-32* 24 -24])^(c[25]&ahead[1023-32* 24 -25])^(c[26]&ahead[1023-32* 24 -26])^(c[27]&ahead[1023-32* 24 -27])^(c[28]&ahead[1023-32* 24 -28])^(c[29]&ahead[1023-32* 24 -29])^(c[30]&ahead[1023-32* 24 -30])^(c[31]&ahead[1023-32* 24 -31]);
  //   newcrc[25]  = (c[0]&ahead[1023-32* 25 ])^(c[1]&ahead[1023-32* 25 -1])^(c[2]&ahead[1023-32* -2 ])^(c[3]&ahead[1023-32* 25 -3])^(c[4]&ahead[1023-32* 25 -4])^(c[5]&ahead[1023-32* 25 -5])^(c[6]&ahead[1023-32* 25 -6])^(c[7]&ahead[1023-32* 25 -7])^(c[8]&ahead[1023-32* 25 -8])^(c[9]&ahead[1023-32* 25 -9])^(c[10]&ahead[1023-32* 25 -10])^(c[11]&ahead[1023-32* 25 -11])^(c[12]&ahead[1023-32* 25 -12])^(c[13]&ahead[1023-32* 25 -13])^(c[14]&ahead[1023-32* 25 -14])^(c[15]&ahead[1023-32* 25 -15])^(c[16]&ahead[1023-32* 25 -16])^(c[17]&ahead[1023-32* 25 -17])^(c[18]&ahead[1023-32* 25 -18])^(c[19]&ahead[1023-32* 25 -19])^(c[20]&ahead[1023-32* 25 -20])^(c[21]&ahead[1023-32* 25 -21])^(c[22]&ahead[1023-32* 25 -22])^(c[23]&ahead[1023-32* 25 -23])^(c[24]&ahead[1023-32* 25 -24])^(c[25]&ahead[1023-32* 25 -25])^(c[26]&ahead[1023-32* 25 -26])^(c[27]&ahead[1023-32* 25 -27])^(c[28]&ahead[1023-32* 25 -28])^(c[29]&ahead[1023-32* 25 -29])^(c[30]&ahead[1023-32* 25 -30])^(c[31]&ahead[1023-32* 25 -31]);
  //   newcrc[26]  = (c[0]&ahead[1023-32* 26 ])^(c[1]&ahead[1023-32* 26 -1])^(c[2]&ahead[1023-32* -2 ])^(c[3]&ahead[1023-32* 26 -3])^(c[4]&ahead[1023-32* 26 -4])^(c[5]&ahead[1023-32* 26 -5])^(c[6]&ahead[1023-32* 26 -6])^(c[7]&ahead[1023-32* 26 -7])^(c[8]&ahead[1023-32* 26 -8])^(c[9]&ahead[1023-32* 26 -9])^(c[10]&ahead[1023-32* 26 -10])^(c[11]&ahead[1023-32* 26 -11])^(c[12]&ahead[1023-32* 26 -12])^(c[13]&ahead[1023-32* 26 -13])^(c[14]&ahead[1023-32* 26 -14])^(c[15]&ahead[1023-32* 26 -15])^(c[16]&ahead[1023-32* 26 -16])^(c[17]&ahead[1023-32* 26 -17])^(c[18]&ahead[1023-32* 26 -18])^(c[19]&ahead[1023-32* 26 -19])^(c[20]&ahead[1023-32* 26 -20])^(c[21]&ahead[1023-32* 26 -21])^(c[22]&ahead[1023-32* 26 -22])^(c[23]&ahead[1023-32* 26 -23])^(c[24]&ahead[1023-32* 26 -24])^(c[25]&ahead[1023-32* 26 -25])^(c[26]&ahead[1023-32* 26 -26])^(c[27]&ahead[1023-32* 26 -27])^(c[28]&ahead[1023-32* 26 -28])^(c[29]&ahead[1023-32* 26 -29])^(c[30]&ahead[1023-32* 26 -30])^(c[31]&ahead[1023-32* 26 -31]);
  //   newcrc[27]  = (c[0]&ahead[1023-32* 27 ])^(c[1]&ahead[1023-32* 27 -1])^(c[2]&ahead[1023-32* -2 ])^(c[3]&ahead[1023-32* 27 -3])^(c[4]&ahead[1023-32* 27 -4])^(c[5]&ahead[1023-32* 27 -5])^(c[6]&ahead[1023-32* 27 -6])^(c[7]&ahead[1023-32* 27 -7])^(c[8]&ahead[1023-32* 27 -8])^(c[9]&ahead[1023-32* 27 -9])^(c[10]&ahead[1023-32* 27 -10])^(c[11]&ahead[1023-32* 27 -11])^(c[12]&ahead[1023-32* 27 -12])^(c[13]&ahead[1023-32* 27 -13])^(c[14]&ahead[1023-32* 27 -14])^(c[15]&ahead[1023-32* 27 -15])^(c[16]&ahead[1023-32* 27 -16])^(c[17]&ahead[1023-32* 27 -17])^(c[18]&ahead[1023-32* 27 -18])^(c[19]&ahead[1023-32* 27 -19])^(c[20]&ahead[1023-32* 27 -20])^(c[21]&ahead[1023-32* 27 -21])^(c[22]&ahead[1023-32* 27 -22])^(c[23]&ahead[1023-32* 27 -23])^(c[24]&ahead[1023-32* 27 -24])^(c[25]&ahead[1023-32* 27 -25])^(c[26]&ahead[1023-32* 27 -26])^(c[27]&ahead[1023-32* 27 -27])^(c[28]&ahead[1023-32* 27 -28])^(c[29]&ahead[1023-32* 27 -29])^(c[30]&ahead[1023-32* 27 -30])^(c[31]&ahead[1023-32* 27 -31]);
  //   newcrc[28]  = (c[0]&ahead[1023-32* 28 ])^(c[1]&ahead[1023-32* 28 -1])^(c[2]&ahead[1023-32* -2 ])^(c[3]&ahead[1023-32* 28 -3])^(c[4]&ahead[1023-32* 28 -4])^(c[5]&ahead[1023-32* 28 -5])^(c[6]&ahead[1023-32* 28 -6])^(c[7]&ahead[1023-32* 28 -7])^(c[8]&ahead[1023-32* 28 -8])^(c[9]&ahead[1023-32* 28 -9])^(c[10]&ahead[1023-32* 28 -10])^(c[11]&ahead[1023-32* 28 -11])^(c[12]&ahead[1023-32* 28 -12])^(c[13]&ahead[1023-32* 28 -13])^(c[14]&ahead[1023-32* 28 -14])^(c[15]&ahead[1023-32* 28 -15])^(c[16]&ahead[1023-32* 28 -16])^(c[17]&ahead[1023-32* 28 -17])^(c[18]&ahead[1023-32* 28 -18])^(c[19]&ahead[1023-32* 28 -19])^(c[20]&ahead[1023-32* 28 -20])^(c[21]&ahead[1023-32* 28 -21])^(c[22]&ahead[1023-32* 28 -22])^(c[23]&ahead[1023-32* 28 -23])^(c[24]&ahead[1023-32* 28 -24])^(c[25]&ahead[1023-32* 28 -25])^(c[26]&ahead[1023-32* 28 -26])^(c[27]&ahead[1023-32* 28 -27])^(c[28]&ahead[1023-32* 28 -28])^(c[29]&ahead[1023-32* 28 -29])^(c[30]&ahead[1023-32* 28 -30])^(c[31]&ahead[1023-32* 28 -31]);
  //   newcrc[29]  = (c[0]&ahead[1023-32* 29 ])^(c[1]&ahead[1023-32* 29 -1])^(c[2]&ahead[1023-32* -2 ])^(c[3]&ahead[1023-32* 29 -3])^(c[4]&ahead[1023-32* 29 -4])^(c[5]&ahead[1023-32* 29 -5])^(c[6]&ahead[1023-32* 29 -6])^(c[7]&ahead[1023-32* 29 -7])^(c[8]&ahead[1023-32* 29 -8])^(c[9]&ahead[1023-32* 29 -9])^(c[10]&ahead[1023-32* 29 -10])^(c[11]&ahead[1023-32* 29 -11])^(c[12]&ahead[1023-32* 29 -12])^(c[13]&ahead[1023-32* 29 -13])^(c[14]&ahead[1023-32* 29 -14])^(c[15]&ahead[1023-32* 29 -15])^(c[16]&ahead[1023-32* 29 -16])^(c[17]&ahead[1023-32* 29 -17])^(c[18]&ahead[1023-32* 29 -18])^(c[19]&ahead[1023-32* 29 -19])^(c[20]&ahead[1023-32* 29 -20])^(c[21]&ahead[1023-32* 29 -21])^(c[22]&ahead[1023-32* 29 -22])^(c[23]&ahead[1023-32* 29 -23])^(c[24]&ahead[1023-32* 29 -24])^(c[25]&ahead[1023-32* 29 -25])^(c[26]&ahead[1023-32* 29 -26])^(c[27]&ahead[1023-32* 29 -27])^(c[28]&ahead[1023-32* 29 -28])^(c[29]&ahead[1023-32* 29 -29])^(c[30]&ahead[1023-32* 29 -30])^(c[31]&ahead[1023-32* 29 -31]);
  //   newcrc[30]  = (c[0]&ahead[1023-32* 30 ])^(c[1]&ahead[1023-32* 30 -1])^(c[2]&ahead[1023-32* -2 ])^(c[3]&ahead[1023-32* 30 -3])^(c[4]&ahead[1023-32* 30 -4])^(c[5]&ahead[1023-32* 30 -5])^(c[6]&ahead[1023-32* 30 -6])^(c[7]&ahead[1023-32* 30 -7])^(c[8]&ahead[1023-32* 30 -8])^(c[9]&ahead[1023-32* 30 -9])^(c[10]&ahead[1023-32* 30 -10])^(c[11]&ahead[1023-32* 30 -11])^(c[12]&ahead[1023-32* 30 -12])^(c[13]&ahead[1023-32* 30 -13])^(c[14]&ahead[1023-32* 30 -14])^(c[15]&ahead[1023-32* 30 -15])^(c[16]&ahead[1023-32* 30 -16])^(c[17]&ahead[1023-32* 30 -17])^(c[18]&ahead[1023-32* 30 -18])^(c[19]&ahead[1023-32* 30 -19])^(c[20]&ahead[1023-32* 30 -20])^(c[21]&ahead[1023-32* 30 -21])^(c[22]&ahead[1023-32* 30 -22])^(c[23]&ahead[1023-32* 30 -23])^(c[24]&ahead[1023-32* 30 -24])^(c[25]&ahead[1023-32* 30 -25])^(c[26]&ahead[1023-32* 30 -26])^(c[27]&ahead[1023-32* 30 -27])^(c[28]&ahead[1023-32* 30 -28])^(c[29]&ahead[1023-32* 30 -29])^(c[30]&ahead[1023-32* 30 -30])^(c[31]&ahead[1023-32* 30 -31]);
  //   newcrc[31]  = (c[0]&ahead[1023-32* 31 ])^(c[1]&ahead[1023-32* 31 -1])^(c[2]&ahead[1023-32* -2 ])^(c[3]&ahead[1023-32* 31 -3])^(c[4]&ahead[1023-32* 31 -4])^(c[5]&ahead[1023-32* 31 -5])^(c[6]&ahead[1023-32* 31 -6])^(c[7]&ahead[1023-32* 31 -7])^(c[8]&ahead[1023-32* 31 -8])^(c[9]&ahead[1023-32* 31 -9])^(c[10]&ahead[1023-32* 31 -10])^(c[11]&ahead[1023-32* 31 -11])^(c[12]&ahead[1023-32* 31 -12])^(c[13]&ahead[1023-32* 31 -13])^(c[14]&ahead[1023-32* 31 -14])^(c[15]&ahead[1023-32* 31 -15])^(c[16]&ahead[1023-32* 31 -16])^(c[17]&ahead[1023-32* 31 -17])^(c[18]&ahead[1023-32* 31 -18])^(c[19]&ahead[1023-32* 31 -19])^(c[20]&ahead[1023-32* 31 -20])^(c[21]&ahead[1023-32* 31 -21])^(c[22]&ahead[1023-32* 31 -22])^(c[23]&ahead[1023-32* 31 -23])^(c[24]&ahead[1023-32* 31 -24])^(c[25]&ahead[1023-32* 31 -25])^(c[26]&ahead[1023-32* 31 -26])^(c[27]&ahead[1023-32* 31 -27])^(c[28]&ahead[1023-32* 31 -28])^(c[29]&ahead[1023-32* 31 -29])^(c[30]&ahead[1023-32* 31 -30])^(c[31]&ahead[1023-32* 31 -31]);
  //   CRC32_ahead = newcrc;
  // end
  // endfunction


// assign test[0 ] =    (crc_i[0]&ahead[1023-32* 0  ])^(crc_i[1]&ahead[1023-32* 0  -1])^(crc_i[2]&ahead[1023-32*0  -2 ])^(crc_i[3]&ahead[1023-32* 0  -3])^(crc_i[4]&ahead[1023-32* 0  -4])^(crc_i[5]&ahead[1023-32* 0  -5])^(crc_i[6]&ahead[1023-32* 0  -6])^(crc_i[7]&ahead[1023-32* 0  -7])^(crc_i[8]&ahead[1023-32* 0  -8])^(crc_i[9]&ahead[1023-32* 0  -9])^(crc_i[10]&ahead[1023-32* 0  -10])^(crc_i[11]&ahead[1023-32* 0  -11])^(crc_i[12]&ahead[1023-32* 0  -12])^(crc_i[13]&ahead[1023-32* 0  -13])^(crc_i[14]&ahead[1023-32* 0  -14])^(crc_i[15]&ahead[1023-32* 0  -15])^(crc_i[16]&ahead[1023-32* 0  -16])^(crc_i[17]&ahead[1023-32* 0  -17])^(crc_i[18]&ahead[1023-32* 0  -18])^(crc_i[19]&ahead[1023-32* 0  -19])^(crc_i[20]&ahead[1023-32* 0  -20])^(crc_i[21]&ahead[1023-32* 0  -21])^(crc_i[22]&ahead[1023-32* 0  -22])^(crc_i[23]&ahead[1023-32* 0  -23])^(crc_i[24]&ahead[1023-32* 0  -24])^(crc_i[25]&ahead[1023-32* 0  -25])^(crc_i[26]&ahead[1023-32* 0  -26])^(crc_i[27]&ahead[1023-32* 0  -27])^(crc_i[28]&ahead[1023-32* 0  -28])^(crc_i[29]&ahead[1023-32* 0  -29])^(crc_i[30]&ahead[1023-32* 0  -30])^(crc_i[31]&ahead[1023-32* 0  -31]);
// assign test[1 ] =    (crc_i[0]&ahead[1023-32* 1  ])^(crc_i[1]&ahead[1023-32* 1  -1])^(crc_i[2]&ahead[1023-32*1  -2 ])^(crc_i[3]&ahead[1023-32* 1  -3])^(crc_i[4]&ahead[1023-32* 1  -4])^(crc_i[5]&ahead[1023-32* 1  -5])^(crc_i[6]&ahead[1023-32* 1  -6])^(crc_i[7]&ahead[1023-32* 1  -7])^(crc_i[8]&ahead[1023-32* 1  -8])^(crc_i[9]&ahead[1023-32* 1  -9])^(crc_i[10]&ahead[1023-32* 1  -10])^(crc_i[11]&ahead[1023-32* 1  -11])^(crc_i[12]&ahead[1023-32* 1  -12])^(crc_i[13]&ahead[1023-32* 1  -13])^(crc_i[14]&ahead[1023-32* 1  -14])^(crc_i[15]&ahead[1023-32* 1  -15])^(crc_i[16]&ahead[1023-32* 1  -16])^(crc_i[17]&ahead[1023-32* 1  -17])^(crc_i[18]&ahead[1023-32* 1  -18])^(crc_i[19]&ahead[1023-32* 1  -19])^(crc_i[20]&ahead[1023-32* 1  -20])^(crc_i[21]&ahead[1023-32* 1  -21])^(crc_i[22]&ahead[1023-32* 1  -22])^(crc_i[23]&ahead[1023-32* 1  -23])^(crc_i[24]&ahead[1023-32* 1  -24])^(crc_i[25]&ahead[1023-32* 1  -25])^(crc_i[26]&ahead[1023-32* 1  -26])^(crc_i[27]&ahead[1023-32* 1  -27])^(crc_i[28]&ahead[1023-32* 1  -28])^(crc_i[29]&ahead[1023-32* 1  -29])^(crc_i[30]&ahead[1023-32* 1  -30])^(crc_i[31]&ahead[1023-32* 1  -31]);
// assign test[2 ] =    (crc_i[0]&ahead[1023-32* 2  ])^(crc_i[1]&ahead[1023-32* 2  -1])^(crc_i[2]&ahead[1023-32*2  -2 ])^(crc_i[3]&ahead[1023-32* 2  -3])^(crc_i[4]&ahead[1023-32* 2  -4])^(crc_i[5]&ahead[1023-32* 2  -5])^(crc_i[6]&ahead[1023-32* 2  -6])^(crc_i[7]&ahead[1023-32* 2  -7])^(crc_i[8]&ahead[1023-32* 2  -8])^(crc_i[9]&ahead[1023-32* 2  -9])^(crc_i[10]&ahead[1023-32* 2  -10])^(crc_i[11]&ahead[1023-32* 2  -11])^(crc_i[12]&ahead[1023-32* 2  -12])^(crc_i[13]&ahead[1023-32* 2  -13])^(crc_i[14]&ahead[1023-32* 2  -14])^(crc_i[15]&ahead[1023-32* 2  -15])^(crc_i[16]&ahead[1023-32* 2  -16])^(crc_i[17]&ahead[1023-32* 2  -17])^(crc_i[18]&ahead[1023-32* 2  -18])^(crc_i[19]&ahead[1023-32* 2  -19])^(crc_i[20]&ahead[1023-32* 2  -20])^(crc_i[21]&ahead[1023-32* 2  -21])^(crc_i[22]&ahead[1023-32* 2  -22])^(crc_i[23]&ahead[1023-32* 2  -23])^(crc_i[24]&ahead[1023-32* 2  -24])^(crc_i[25]&ahead[1023-32* 2  -25])^(crc_i[26]&ahead[1023-32* 2  -26])^(crc_i[27]&ahead[1023-32* 2  -27])^(crc_i[28]&ahead[1023-32* 2  -28])^(crc_i[29]&ahead[1023-32* 2  -29])^(crc_i[30]&ahead[1023-32* 2  -30])^(crc_i[31]&ahead[1023-32* 2  -31]);
// assign test[3 ] =    (crc_i[0]&ahead[1023-32* 3  ])^(crc_i[1]&ahead[1023-32* 3  -1])^(crc_i[2]&ahead[1023-32*3  -2 ])^(crc_i[3]&ahead[1023-32* 3  -3])^(crc_i[4]&ahead[1023-32* 3  -4])^(crc_i[5]&ahead[1023-32* 3  -5])^(crc_i[6]&ahead[1023-32* 3  -6])^(crc_i[7]&ahead[1023-32* 3  -7])^(crc_i[8]&ahead[1023-32* 3  -8])^(crc_i[9]&ahead[1023-32* 3  -9])^(crc_i[10]&ahead[1023-32* 3  -10])^(crc_i[11]&ahead[1023-32* 3  -11])^(crc_i[12]&ahead[1023-32* 3  -12])^(crc_i[13]&ahead[1023-32* 3  -13])^(crc_i[14]&ahead[1023-32* 3  -14])^(crc_i[15]&ahead[1023-32* 3  -15])^(crc_i[16]&ahead[1023-32* 3  -16])^(crc_i[17]&ahead[1023-32* 3  -17])^(crc_i[18]&ahead[1023-32* 3  -18])^(crc_i[19]&ahead[1023-32* 3  -19])^(crc_i[20]&ahead[1023-32* 3  -20])^(crc_i[21]&ahead[1023-32* 3  -21])^(crc_i[22]&ahead[1023-32* 3  -22])^(crc_i[23]&ahead[1023-32* 3  -23])^(crc_i[24]&ahead[1023-32* 3  -24])^(crc_i[25]&ahead[1023-32* 3  -25])^(crc_i[26]&ahead[1023-32* 3  -26])^(crc_i[27]&ahead[1023-32* 3  -27])^(crc_i[28]&ahead[1023-32* 3  -28])^(crc_i[29]&ahead[1023-32* 3  -29])^(crc_i[30]&ahead[1023-32* 3  -30])^(crc_i[31]&ahead[1023-32* 3  -31]);
// assign test[4 ] =    (crc_i[0]&ahead[1023-32* 4  ])^(crc_i[1]&ahead[1023-32* 4  -1])^(crc_i[2]&ahead[1023-32*4  -2 ])^(crc_i[3]&ahead[1023-32* 4  -3])^(crc_i[4]&ahead[1023-32* 4  -4])^(crc_i[5]&ahead[1023-32* 4  -5])^(crc_i[6]&ahead[1023-32* 4  -6])^(crc_i[7]&ahead[1023-32* 4  -7])^(crc_i[8]&ahead[1023-32* 4  -8])^(crc_i[9]&ahead[1023-32* 4  -9])^(crc_i[10]&ahead[1023-32* 4  -10])^(crc_i[11]&ahead[1023-32* 4  -11])^(crc_i[12]&ahead[1023-32* 4  -12])^(crc_i[13]&ahead[1023-32* 4  -13])^(crc_i[14]&ahead[1023-32* 4  -14])^(crc_i[15]&ahead[1023-32* 4  -15])^(crc_i[16]&ahead[1023-32* 4  -16])^(crc_i[17]&ahead[1023-32* 4  -17])^(crc_i[18]&ahead[1023-32* 4  -18])^(crc_i[19]&ahead[1023-32* 4  -19])^(crc_i[20]&ahead[1023-32* 4  -20])^(crc_i[21]&ahead[1023-32* 4  -21])^(crc_i[22]&ahead[1023-32* 4  -22])^(crc_i[23]&ahead[1023-32* 4  -23])^(crc_i[24]&ahead[1023-32* 4  -24])^(crc_i[25]&ahead[1023-32* 4  -25])^(crc_i[26]&ahead[1023-32* 4  -26])^(crc_i[27]&ahead[1023-32* 4  -27])^(crc_i[28]&ahead[1023-32* 4  -28])^(crc_i[29]&ahead[1023-32* 4  -29])^(crc_i[30]&ahead[1023-32* 4  -30])^(crc_i[31]&ahead[1023-32* 4  -31]);
// assign test[5 ] =    (crc_i[0]&ahead[1023-32* 5  ])^(crc_i[1]&ahead[1023-32* 5  -1])^(crc_i[2]&ahead[1023-32*5  -2 ])^(crc_i[3]&ahead[1023-32* 5  -3])^(crc_i[4]&ahead[1023-32* 5  -4])^(crc_i[5]&ahead[1023-32* 5  -5])^(crc_i[6]&ahead[1023-32* 5  -6])^(crc_i[7]&ahead[1023-32* 5  -7])^(crc_i[8]&ahead[1023-32* 5  -8])^(crc_i[9]&ahead[1023-32* 5  -9])^(crc_i[10]&ahead[1023-32* 5  -10])^(crc_i[11]&ahead[1023-32* 5  -11])^(crc_i[12]&ahead[1023-32* 5  -12])^(crc_i[13]&ahead[1023-32* 5  -13])^(crc_i[14]&ahead[1023-32* 5  -14])^(crc_i[15]&ahead[1023-32* 5  -15])^(crc_i[16]&ahead[1023-32* 5  -16])^(crc_i[17]&ahead[1023-32* 5  -17])^(crc_i[18]&ahead[1023-32* 5  -18])^(crc_i[19]&ahead[1023-32* 5  -19])^(crc_i[20]&ahead[1023-32* 5  -20])^(crc_i[21]&ahead[1023-32* 5  -21])^(crc_i[22]&ahead[1023-32* 5  -22])^(crc_i[23]&ahead[1023-32* 5  -23])^(crc_i[24]&ahead[1023-32* 5  -24])^(crc_i[25]&ahead[1023-32* 5  -25])^(crc_i[26]&ahead[1023-32* 5  -26])^(crc_i[27]&ahead[1023-32* 5  -27])^(crc_i[28]&ahead[1023-32* 5  -28])^(crc_i[29]&ahead[1023-32* 5  -29])^(crc_i[30]&ahead[1023-32* 5  -30])^(crc_i[31]&ahead[1023-32* 5  -31]);
// assign test[6 ] =    (crc_i[0]&ahead[1023-32* 6  ])^(crc_i[1]&ahead[1023-32* 6  -1])^(crc_i[2]&ahead[1023-32*6  -2 ])^(crc_i[3]&ahead[1023-32* 6  -3])^(crc_i[4]&ahead[1023-32* 6  -4])^(crc_i[5]&ahead[1023-32* 6  -5])^(crc_i[6]&ahead[1023-32* 6  -6])^(crc_i[7]&ahead[1023-32* 6  -7])^(crc_i[8]&ahead[1023-32* 6  -8])^(crc_i[9]&ahead[1023-32* 6  -9])^(crc_i[10]&ahead[1023-32* 6  -10])^(crc_i[11]&ahead[1023-32* 6  -11])^(crc_i[12]&ahead[1023-32* 6  -12])^(crc_i[13]&ahead[1023-32* 6  -13])^(crc_i[14]&ahead[1023-32* 6  -14])^(crc_i[15]&ahead[1023-32* 6  -15])^(crc_i[16]&ahead[1023-32* 6  -16])^(crc_i[17]&ahead[1023-32* 6  -17])^(crc_i[18]&ahead[1023-32* 6  -18])^(crc_i[19]&ahead[1023-32* 6  -19])^(crc_i[20]&ahead[1023-32* 6  -20])^(crc_i[21]&ahead[1023-32* 6  -21])^(crc_i[22]&ahead[1023-32* 6  -22])^(crc_i[23]&ahead[1023-32* 6  -23])^(crc_i[24]&ahead[1023-32* 6  -24])^(crc_i[25]&ahead[1023-32* 6  -25])^(crc_i[26]&ahead[1023-32* 6  -26])^(crc_i[27]&ahead[1023-32* 6  -27])^(crc_i[28]&ahead[1023-32* 6  -28])^(crc_i[29]&ahead[1023-32* 6  -29])^(crc_i[30]&ahead[1023-32* 6  -30])^(crc_i[31]&ahead[1023-32* 6  -31]);
// assign test[7 ] =    (crc_i[0]&ahead[1023-32* 7  ])^(crc_i[1]&ahead[1023-32* 7  -1])^(crc_i[2]&ahead[1023-32*7  -2 ])^(crc_i[3]&ahead[1023-32* 7  -3])^(crc_i[4]&ahead[1023-32* 7  -4])^(crc_i[5]&ahead[1023-32* 7  -5])^(crc_i[6]&ahead[1023-32* 7  -6])^(crc_i[7]&ahead[1023-32* 7  -7])^(crc_i[8]&ahead[1023-32* 7  -8])^(crc_i[9]&ahead[1023-32* 7  -9])^(crc_i[10]&ahead[1023-32* 7  -10])^(crc_i[11]&ahead[1023-32* 7  -11])^(crc_i[12]&ahead[1023-32* 7  -12])^(crc_i[13]&ahead[1023-32* 7  -13])^(crc_i[14]&ahead[1023-32* 7  -14])^(crc_i[15]&ahead[1023-32* 7  -15])^(crc_i[16]&ahead[1023-32* 7  -16])^(crc_i[17]&ahead[1023-32* 7  -17])^(crc_i[18]&ahead[1023-32* 7  -18])^(crc_i[19]&ahead[1023-32* 7  -19])^(crc_i[20]&ahead[1023-32* 7  -20])^(crc_i[21]&ahead[1023-32* 7  -21])^(crc_i[22]&ahead[1023-32* 7  -22])^(crc_i[23]&ahead[1023-32* 7  -23])^(crc_i[24]&ahead[1023-32* 7  -24])^(crc_i[25]&ahead[1023-32* 7  -25])^(crc_i[26]&ahead[1023-32* 7  -26])^(crc_i[27]&ahead[1023-32* 7  -27])^(crc_i[28]&ahead[1023-32* 7  -28])^(crc_i[29]&ahead[1023-32* 7  -29])^(crc_i[30]&ahead[1023-32* 7  -30])^(crc_i[31]&ahead[1023-32* 7  -31]);
// assign test[8 ] =    (crc_i[0]&ahead[1023-32* 8  ])^(crc_i[1]&ahead[1023-32* 8  -1])^(crc_i[2]&ahead[1023-32*8  -2 ])^(crc_i[3]&ahead[1023-32* 8  -3])^(crc_i[4]&ahead[1023-32* 8  -4])^(crc_i[5]&ahead[1023-32* 8  -5])^(crc_i[6]&ahead[1023-32* 8  -6])^(crc_i[7]&ahead[1023-32* 8  -7])^(crc_i[8]&ahead[1023-32* 8  -8])^(crc_i[9]&ahead[1023-32* 8  -9])^(crc_i[10]&ahead[1023-32* 8  -10])^(crc_i[11]&ahead[1023-32* 8  -11])^(crc_i[12]&ahead[1023-32* 8  -12])^(crc_i[13]&ahead[1023-32* 8  -13])^(crc_i[14]&ahead[1023-32* 8  -14])^(crc_i[15]&ahead[1023-32* 8  -15])^(crc_i[16]&ahead[1023-32* 8  -16])^(crc_i[17]&ahead[1023-32* 8  -17])^(crc_i[18]&ahead[1023-32* 8  -18])^(crc_i[19]&ahead[1023-32* 8  -19])^(crc_i[20]&ahead[1023-32* 8  -20])^(crc_i[21]&ahead[1023-32* 8  -21])^(crc_i[22]&ahead[1023-32* 8  -22])^(crc_i[23]&ahead[1023-32* 8  -23])^(crc_i[24]&ahead[1023-32* 8  -24])^(crc_i[25]&ahead[1023-32* 8  -25])^(crc_i[26]&ahead[1023-32* 8  -26])^(crc_i[27]&ahead[1023-32* 8  -27])^(crc_i[28]&ahead[1023-32* 8  -28])^(crc_i[29]&ahead[1023-32* 8  -29])^(crc_i[30]&ahead[1023-32* 8  -30])^(crc_i[31]&ahead[1023-32* 8  -31]);
// assign test[9 ] =    (crc_i[0]&ahead[1023-32* 9  ])^(crc_i[1]&ahead[1023-32* 9  -1])^(crc_i[2]&ahead[1023-32*9  -2 ])^(crc_i[3]&ahead[1023-32* 9  -3])^(crc_i[4]&ahead[1023-32* 9  -4])^(crc_i[5]&ahead[1023-32* 9  -5])^(crc_i[6]&ahead[1023-32* 9  -6])^(crc_i[7]&ahead[1023-32* 9  -7])^(crc_i[8]&ahead[1023-32* 9  -8])^(crc_i[9]&ahead[1023-32* 9  -9])^(crc_i[10]&ahead[1023-32* 9  -10])^(crc_i[11]&ahead[1023-32* 9  -11])^(crc_i[12]&ahead[1023-32* 9  -12])^(crc_i[13]&ahead[1023-32* 9  -13])^(crc_i[14]&ahead[1023-32* 9  -14])^(crc_i[15]&ahead[1023-32* 9  -15])^(crc_i[16]&ahead[1023-32* 9  -16])^(crc_i[17]&ahead[1023-32* 9  -17])^(crc_i[18]&ahead[1023-32* 9  -18])^(crc_i[19]&ahead[1023-32* 9  -19])^(crc_i[20]&ahead[1023-32* 9  -20])^(crc_i[21]&ahead[1023-32* 9  -21])^(crc_i[22]&ahead[1023-32* 9  -22])^(crc_i[23]&ahead[1023-32* 9  -23])^(crc_i[24]&ahead[1023-32* 9  -24])^(crc_i[25]&ahead[1023-32* 9  -25])^(crc_i[26]&ahead[1023-32* 9  -26])^(crc_i[27]&ahead[1023-32* 9  -27])^(crc_i[28]&ahead[1023-32* 9  -28])^(crc_i[29]&ahead[1023-32* 9  -29])^(crc_i[30]&ahead[1023-32* 9  -30])^(crc_i[31]&ahead[1023-32* 9  -31]);
// assign test[10] =    (crc_i[0]&ahead[1023-32* 10 ])^(crc_i[1]&ahead[1023-32* 10 -1])^(crc_i[2]&ahead[1023-32*10 -2 ])^(crc_i[3]&ahead[1023-32* 10 -3])^(crc_i[4]&ahead[1023-32* 10 -4])^(crc_i[5]&ahead[1023-32* 10 -5])^(crc_i[6]&ahead[1023-32* 10 -6])^(crc_i[7]&ahead[1023-32* 10 -7])^(crc_i[8]&ahead[1023-32* 10 -8])^(crc_i[9]&ahead[1023-32* 10 -9])^(crc_i[10]&ahead[1023-32* 10 -10])^(crc_i[11]&ahead[1023-32* 10 -11])^(crc_i[12]&ahead[1023-32* 10 -12])^(crc_i[13]&ahead[1023-32* 10 -13])^(crc_i[14]&ahead[1023-32* 10 -14])^(crc_i[15]&ahead[1023-32* 10 -15])^(crc_i[16]&ahead[1023-32* 10 -16])^(crc_i[17]&ahead[1023-32* 10 -17])^(crc_i[18]&ahead[1023-32* 10 -18])^(crc_i[19]&ahead[1023-32* 10 -19])^(crc_i[20]&ahead[1023-32* 10 -20])^(crc_i[21]&ahead[1023-32* 10 -21])^(crc_i[22]&ahead[1023-32* 10 -22])^(crc_i[23]&ahead[1023-32* 10 -23])^(crc_i[24]&ahead[1023-32* 10 -24])^(crc_i[25]&ahead[1023-32* 10 -25])^(crc_i[26]&ahead[1023-32* 10 -26])^(crc_i[27]&ahead[1023-32* 10 -27])^(crc_i[28]&ahead[1023-32* 10 -28])^(crc_i[29]&ahead[1023-32* 10 -29])^(crc_i[30]&ahead[1023-32* 10 -30])^(crc_i[31]&ahead[1023-32* 10 -31]);
// assign test[11] =    (crc_i[0]&ahead[1023-32* 11 ])^(crc_i[1]&ahead[1023-32* 11 -1])^(crc_i[2]&ahead[1023-32*11 -2 ])^(crc_i[3]&ahead[1023-32* 11 -3])^(crc_i[4]&ahead[1023-32* 11 -4])^(crc_i[5]&ahead[1023-32* 11 -5])^(crc_i[6]&ahead[1023-32* 11 -6])^(crc_i[7]&ahead[1023-32* 11 -7])^(crc_i[8]&ahead[1023-32* 11 -8])^(crc_i[9]&ahead[1023-32* 11 -9])^(crc_i[10]&ahead[1023-32* 11 -10])^(crc_i[11]&ahead[1023-32* 11 -11])^(crc_i[12]&ahead[1023-32* 11 -12])^(crc_i[13]&ahead[1023-32* 11 -13])^(crc_i[14]&ahead[1023-32* 11 -14])^(crc_i[15]&ahead[1023-32* 11 -15])^(crc_i[16]&ahead[1023-32* 11 -16])^(crc_i[17]&ahead[1023-32* 11 -17])^(crc_i[18]&ahead[1023-32* 11 -18])^(crc_i[19]&ahead[1023-32* 11 -19])^(crc_i[20]&ahead[1023-32* 11 -20])^(crc_i[21]&ahead[1023-32* 11 -21])^(crc_i[22]&ahead[1023-32* 11 -22])^(crc_i[23]&ahead[1023-32* 11 -23])^(crc_i[24]&ahead[1023-32* 11 -24])^(crc_i[25]&ahead[1023-32* 11 -25])^(crc_i[26]&ahead[1023-32* 11 -26])^(crc_i[27]&ahead[1023-32* 11 -27])^(crc_i[28]&ahead[1023-32* 11 -28])^(crc_i[29]&ahead[1023-32* 11 -29])^(crc_i[30]&ahead[1023-32* 11 -30])^(crc_i[31]&ahead[1023-32* 11 -31]);
// assign test[12] =    (crc_i[0]&ahead[1023-32* 12 ])^(crc_i[1]&ahead[1023-32* 12 -1])^(crc_i[2]&ahead[1023-32*12 -2 ])^(crc_i[3]&ahead[1023-32* 12 -3])^(crc_i[4]&ahead[1023-32* 12 -4])^(crc_i[5]&ahead[1023-32* 12 -5])^(crc_i[6]&ahead[1023-32* 12 -6])^(crc_i[7]&ahead[1023-32* 12 -7])^(crc_i[8]&ahead[1023-32* 12 -8])^(crc_i[9]&ahead[1023-32* 12 -9])^(crc_i[10]&ahead[1023-32* 12 -10])^(crc_i[11]&ahead[1023-32* 12 -11])^(crc_i[12]&ahead[1023-32* 12 -12])^(crc_i[13]&ahead[1023-32* 12 -13])^(crc_i[14]&ahead[1023-32* 12 -14])^(crc_i[15]&ahead[1023-32* 12 -15])^(crc_i[16]&ahead[1023-32* 12 -16])^(crc_i[17]&ahead[1023-32* 12 -17])^(crc_i[18]&ahead[1023-32* 12 -18])^(crc_i[19]&ahead[1023-32* 12 -19])^(crc_i[20]&ahead[1023-32* 12 -20])^(crc_i[21]&ahead[1023-32* 12 -21])^(crc_i[22]&ahead[1023-32* 12 -22])^(crc_i[23]&ahead[1023-32* 12 -23])^(crc_i[24]&ahead[1023-32* 12 -24])^(crc_i[25]&ahead[1023-32* 12 -25])^(crc_i[26]&ahead[1023-32* 12 -26])^(crc_i[27]&ahead[1023-32* 12 -27])^(crc_i[28]&ahead[1023-32* 12 -28])^(crc_i[29]&ahead[1023-32* 12 -29])^(crc_i[30]&ahead[1023-32* 12 -30])^(crc_i[31]&ahead[1023-32* 12 -31]);
// assign test[13] =    (crc_i[0]&ahead[1023-32* 13 ])^(crc_i[1]&ahead[1023-32* 13 -1])^(crc_i[2]&ahead[1023-32*13 -2 ])^(crc_i[3]&ahead[1023-32* 13 -3])^(crc_i[4]&ahead[1023-32* 13 -4])^(crc_i[5]&ahead[1023-32* 13 -5])^(crc_i[6]&ahead[1023-32* 13 -6])^(crc_i[7]&ahead[1023-32* 13 -7])^(crc_i[8]&ahead[1023-32* 13 -8])^(crc_i[9]&ahead[1023-32* 13 -9])^(crc_i[10]&ahead[1023-32* 13 -10])^(crc_i[11]&ahead[1023-32* 13 -11])^(crc_i[12]&ahead[1023-32* 13 -12])^(crc_i[13]&ahead[1023-32* 13 -13])^(crc_i[14]&ahead[1023-32* 13 -14])^(crc_i[15]&ahead[1023-32* 13 -15])^(crc_i[16]&ahead[1023-32* 13 -16])^(crc_i[17]&ahead[1023-32* 13 -17])^(crc_i[18]&ahead[1023-32* 13 -18])^(crc_i[19]&ahead[1023-32* 13 -19])^(crc_i[20]&ahead[1023-32* 13 -20])^(crc_i[21]&ahead[1023-32* 13 -21])^(crc_i[22]&ahead[1023-32* 13 -22])^(crc_i[23]&ahead[1023-32* 13 -23])^(crc_i[24]&ahead[1023-32* 13 -24])^(crc_i[25]&ahead[1023-32* 13 -25])^(crc_i[26]&ahead[1023-32* 13 -26])^(crc_i[27]&ahead[1023-32* 13 -27])^(crc_i[28]&ahead[1023-32* 13 -28])^(crc_i[29]&ahead[1023-32* 13 -29])^(crc_i[30]&ahead[1023-32* 13 -30])^(crc_i[31]&ahead[1023-32* 13 -31]);
// assign test[14] =    (crc_i[0]&ahead[1023-32* 14 ])^(crc_i[1]&ahead[1023-32* 14 -1])^(crc_i[2]&ahead[1023-32*14 -2 ])^(crc_i[3]&ahead[1023-32* 14 -3])^(crc_i[4]&ahead[1023-32* 14 -4])^(crc_i[5]&ahead[1023-32* 14 -5])^(crc_i[6]&ahead[1023-32* 14 -6])^(crc_i[7]&ahead[1023-32* 14 -7])^(crc_i[8]&ahead[1023-32* 14 -8])^(crc_i[9]&ahead[1023-32* 14 -9])^(crc_i[10]&ahead[1023-32* 14 -10])^(crc_i[11]&ahead[1023-32* 14 -11])^(crc_i[12]&ahead[1023-32* 14 -12])^(crc_i[13]&ahead[1023-32* 14 -13])^(crc_i[14]&ahead[1023-32* 14 -14])^(crc_i[15]&ahead[1023-32* 14 -15])^(crc_i[16]&ahead[1023-32* 14 -16])^(crc_i[17]&ahead[1023-32* 14 -17])^(crc_i[18]&ahead[1023-32* 14 -18])^(crc_i[19]&ahead[1023-32* 14 -19])^(crc_i[20]&ahead[1023-32* 14 -20])^(crc_i[21]&ahead[1023-32* 14 -21])^(crc_i[22]&ahead[1023-32* 14 -22])^(crc_i[23]&ahead[1023-32* 14 -23])^(crc_i[24]&ahead[1023-32* 14 -24])^(crc_i[25]&ahead[1023-32* 14 -25])^(crc_i[26]&ahead[1023-32* 14 -26])^(crc_i[27]&ahead[1023-32* 14 -27])^(crc_i[28]&ahead[1023-32* 14 -28])^(crc_i[29]&ahead[1023-32* 14 -29])^(crc_i[30]&ahead[1023-32* 14 -30])^(crc_i[31]&ahead[1023-32* 14 -31]);
// assign test[15] =    (crc_i[0]&ahead[1023-32* 15 ])^(crc_i[1]&ahead[1023-32* 15 -1])^(crc_i[2]&ahead[1023-32*15 -2 ])^(crc_i[3]&ahead[1023-32* 15 -3])^(crc_i[4]&ahead[1023-32* 15 -4])^(crc_i[5]&ahead[1023-32* 15 -5])^(crc_i[6]&ahead[1023-32* 15 -6])^(crc_i[7]&ahead[1023-32* 15 -7])^(crc_i[8]&ahead[1023-32* 15 -8])^(crc_i[9]&ahead[1023-32* 15 -9])^(crc_i[10]&ahead[1023-32* 15 -10])^(crc_i[11]&ahead[1023-32* 15 -11])^(crc_i[12]&ahead[1023-32* 15 -12])^(crc_i[13]&ahead[1023-32* 15 -13])^(crc_i[14]&ahead[1023-32* 15 -14])^(crc_i[15]&ahead[1023-32* 15 -15])^(crc_i[16]&ahead[1023-32* 15 -16])^(crc_i[17]&ahead[1023-32* 15 -17])^(crc_i[18]&ahead[1023-32* 15 -18])^(crc_i[19]&ahead[1023-32* 15 -19])^(crc_i[20]&ahead[1023-32* 15 -20])^(crc_i[21]&ahead[1023-32* 15 -21])^(crc_i[22]&ahead[1023-32* 15 -22])^(crc_i[23]&ahead[1023-32* 15 -23])^(crc_i[24]&ahead[1023-32* 15 -24])^(crc_i[25]&ahead[1023-32* 15 -25])^(crc_i[26]&ahead[1023-32* 15 -26])^(crc_i[27]&ahead[1023-32* 15 -27])^(crc_i[28]&ahead[1023-32* 15 -28])^(crc_i[29]&ahead[1023-32* 15 -29])^(crc_i[30]&ahead[1023-32* 15 -30])^(crc_i[31]&ahead[1023-32* 15 -31]);
// assign test[16] =    (crc_i[0]&ahead[1023-32* 16 ])^(crc_i[1]&ahead[1023-32* 16 -1])^(crc_i[2]&ahead[1023-32*16 -2 ])^(crc_i[3]&ahead[1023-32* 16 -3])^(crc_i[4]&ahead[1023-32* 16 -4])^(crc_i[5]&ahead[1023-32* 16 -5])^(crc_i[6]&ahead[1023-32* 16 -6])^(crc_i[7]&ahead[1023-32* 16 -7])^(crc_i[8]&ahead[1023-32* 16 -8])^(crc_i[9]&ahead[1023-32* 16 -9])^(crc_i[10]&ahead[1023-32* 16 -10])^(crc_i[11]&ahead[1023-32* 16 -11])^(crc_i[12]&ahead[1023-32* 16 -12])^(crc_i[13]&ahead[1023-32* 16 -13])^(crc_i[14]&ahead[1023-32* 16 -14])^(crc_i[15]&ahead[1023-32* 16 -15])^(crc_i[16]&ahead[1023-32* 16 -16])^(crc_i[17]&ahead[1023-32* 16 -17])^(crc_i[18]&ahead[1023-32* 16 -18])^(crc_i[19]&ahead[1023-32* 16 -19])^(crc_i[20]&ahead[1023-32* 16 -20])^(crc_i[21]&ahead[1023-32* 16 -21])^(crc_i[22]&ahead[1023-32* 16 -22])^(crc_i[23]&ahead[1023-32* 16 -23])^(crc_i[24]&ahead[1023-32* 16 -24])^(crc_i[25]&ahead[1023-32* 16 -25])^(crc_i[26]&ahead[1023-32* 16 -26])^(crc_i[27]&ahead[1023-32* 16 -27])^(crc_i[28]&ahead[1023-32* 16 -28])^(crc_i[29]&ahead[1023-32* 16 -29])^(crc_i[30]&ahead[1023-32* 16 -30])^(crc_i[31]&ahead[1023-32* 16 -31]);
// assign test[17] =    (crc_i[0]&ahead[1023-32* 17 ])^(crc_i[1]&ahead[1023-32* 17 -1])^(crc_i[2]&ahead[1023-32*17 -2 ])^(crc_i[3]&ahead[1023-32* 17 -3])^(crc_i[4]&ahead[1023-32* 17 -4])^(crc_i[5]&ahead[1023-32* 17 -5])^(crc_i[6]&ahead[1023-32* 17 -6])^(crc_i[7]&ahead[1023-32* 17 -7])^(crc_i[8]&ahead[1023-32* 17 -8])^(crc_i[9]&ahead[1023-32* 17 -9])^(crc_i[10]&ahead[1023-32* 17 -10])^(crc_i[11]&ahead[1023-32* 17 -11])^(crc_i[12]&ahead[1023-32* 17 -12])^(crc_i[13]&ahead[1023-32* 17 -13])^(crc_i[14]&ahead[1023-32* 17 -14])^(crc_i[15]&ahead[1023-32* 17 -15])^(crc_i[16]&ahead[1023-32* 17 -16])^(crc_i[17]&ahead[1023-32* 17 -17])^(crc_i[18]&ahead[1023-32* 17 -18])^(crc_i[19]&ahead[1023-32* 17 -19])^(crc_i[20]&ahead[1023-32* 17 -20])^(crc_i[21]&ahead[1023-32* 17 -21])^(crc_i[22]&ahead[1023-32* 17 -22])^(crc_i[23]&ahead[1023-32* 17 -23])^(crc_i[24]&ahead[1023-32* 17 -24])^(crc_i[25]&ahead[1023-32* 17 -25])^(crc_i[26]&ahead[1023-32* 17 -26])^(crc_i[27]&ahead[1023-32* 17 -27])^(crc_i[28]&ahead[1023-32* 17 -28])^(crc_i[29]&ahead[1023-32* 17 -29])^(crc_i[30]&ahead[1023-32* 17 -30])^(crc_i[31]&ahead[1023-32* 17 -31]);
// assign test[18] =    (crc_i[0]&ahead[1023-32* 18 ])^(crc_i[1]&ahead[1023-32* 18 -1])^(crc_i[2]&ahead[1023-32*18 -2 ])^(crc_i[3]&ahead[1023-32* 18 -3])^(crc_i[4]&ahead[1023-32* 18 -4])^(crc_i[5]&ahead[1023-32* 18 -5])^(crc_i[6]&ahead[1023-32* 18 -6])^(crc_i[7]&ahead[1023-32* 18 -7])^(crc_i[8]&ahead[1023-32* 18 -8])^(crc_i[9]&ahead[1023-32* 18 -9])^(crc_i[10]&ahead[1023-32* 18 -10])^(crc_i[11]&ahead[1023-32* 18 -11])^(crc_i[12]&ahead[1023-32* 18 -12])^(crc_i[13]&ahead[1023-32* 18 -13])^(crc_i[14]&ahead[1023-32* 18 -14])^(crc_i[15]&ahead[1023-32* 18 -15])^(crc_i[16]&ahead[1023-32* 18 -16])^(crc_i[17]&ahead[1023-32* 18 -17])^(crc_i[18]&ahead[1023-32* 18 -18])^(crc_i[19]&ahead[1023-32* 18 -19])^(crc_i[20]&ahead[1023-32* 18 -20])^(crc_i[21]&ahead[1023-32* 18 -21])^(crc_i[22]&ahead[1023-32* 18 -22])^(crc_i[23]&ahead[1023-32* 18 -23])^(crc_i[24]&ahead[1023-32* 18 -24])^(crc_i[25]&ahead[1023-32* 18 -25])^(crc_i[26]&ahead[1023-32* 18 -26])^(crc_i[27]&ahead[1023-32* 18 -27])^(crc_i[28]&ahead[1023-32* 18 -28])^(crc_i[29]&ahead[1023-32* 18 -29])^(crc_i[30]&ahead[1023-32* 18 -30])^(crc_i[31]&ahead[1023-32* 18 -31]);
// assign test[19] =    (crc_i[0]&ahead[1023-32* 19 ])^(crc_i[1]&ahead[1023-32* 19 -1])^(crc_i[2]&ahead[1023-32*19 -2 ])^(crc_i[3]&ahead[1023-32* 19 -3])^(crc_i[4]&ahead[1023-32* 19 -4])^(crc_i[5]&ahead[1023-32* 19 -5])^(crc_i[6]&ahead[1023-32* 19 -6])^(crc_i[7]&ahead[1023-32* 19 -7])^(crc_i[8]&ahead[1023-32* 19 -8])^(crc_i[9]&ahead[1023-32* 19 -9])^(crc_i[10]&ahead[1023-32* 19 -10])^(crc_i[11]&ahead[1023-32* 19 -11])^(crc_i[12]&ahead[1023-32* 19 -12])^(crc_i[13]&ahead[1023-32* 19 -13])^(crc_i[14]&ahead[1023-32* 19 -14])^(crc_i[15]&ahead[1023-32* 19 -15])^(crc_i[16]&ahead[1023-32* 19 -16])^(crc_i[17]&ahead[1023-32* 19 -17])^(crc_i[18]&ahead[1023-32* 19 -18])^(crc_i[19]&ahead[1023-32* 19 -19])^(crc_i[20]&ahead[1023-32* 19 -20])^(crc_i[21]&ahead[1023-32* 19 -21])^(crc_i[22]&ahead[1023-32* 19 -22])^(crc_i[23]&ahead[1023-32* 19 -23])^(crc_i[24]&ahead[1023-32* 19 -24])^(crc_i[25]&ahead[1023-32* 19 -25])^(crc_i[26]&ahead[1023-32* 19 -26])^(crc_i[27]&ahead[1023-32* 19 -27])^(crc_i[28]&ahead[1023-32* 19 -28])^(crc_i[29]&ahead[1023-32* 19 -29])^(crc_i[30]&ahead[1023-32* 19 -30])^(crc_i[31]&ahead[1023-32* 19 -31]);
// assign test[20] =    (crc_i[0]&ahead[1023-32* 20 ])^(crc_i[1]&ahead[1023-32* 20 -1])^(crc_i[2]&ahead[1023-32*20 -2 ])^(crc_i[3]&ahead[1023-32* 20 -3])^(crc_i[4]&ahead[1023-32* 20 -4])^(crc_i[5]&ahead[1023-32* 20 -5])^(crc_i[6]&ahead[1023-32* 20 -6])^(crc_i[7]&ahead[1023-32* 20 -7])^(crc_i[8]&ahead[1023-32* 20 -8])^(crc_i[9]&ahead[1023-32* 20 -9])^(crc_i[10]&ahead[1023-32* 20 -10])^(crc_i[11]&ahead[1023-32* 20 -11])^(crc_i[12]&ahead[1023-32* 20 -12])^(crc_i[13]&ahead[1023-32* 20 -13])^(crc_i[14]&ahead[1023-32* 20 -14])^(crc_i[15]&ahead[1023-32* 20 -15])^(crc_i[16]&ahead[1023-32* 20 -16])^(crc_i[17]&ahead[1023-32* 20 -17])^(crc_i[18]&ahead[1023-32* 20 -18])^(crc_i[19]&ahead[1023-32* 20 -19])^(crc_i[20]&ahead[1023-32* 20 -20])^(crc_i[21]&ahead[1023-32* 20 -21])^(crc_i[22]&ahead[1023-32* 20 -22])^(crc_i[23]&ahead[1023-32* 20 -23])^(crc_i[24]&ahead[1023-32* 20 -24])^(crc_i[25]&ahead[1023-32* 20 -25])^(crc_i[26]&ahead[1023-32* 20 -26])^(crc_i[27]&ahead[1023-32* 20 -27])^(crc_i[28]&ahead[1023-32* 20 -28])^(crc_i[29]&ahead[1023-32* 20 -29])^(crc_i[30]&ahead[1023-32* 20 -30])^(crc_i[31]&ahead[1023-32* 20 -31]);
// assign test[21] =    (crc_i[0]&ahead[1023-32* 21 ])^(crc_i[1]&ahead[1023-32* 21 -1])^(crc_i[2]&ahead[1023-32*21 -2 ])^(crc_i[3]&ahead[1023-32* 21 -3])^(crc_i[4]&ahead[1023-32* 21 -4])^(crc_i[5]&ahead[1023-32* 21 -5])^(crc_i[6]&ahead[1023-32* 21 -6])^(crc_i[7]&ahead[1023-32* 21 -7])^(crc_i[8]&ahead[1023-32* 21 -8])^(crc_i[9]&ahead[1023-32* 21 -9])^(crc_i[10]&ahead[1023-32* 21 -10])^(crc_i[11]&ahead[1023-32* 21 -11])^(crc_i[12]&ahead[1023-32* 21 -12])^(crc_i[13]&ahead[1023-32* 21 -13])^(crc_i[14]&ahead[1023-32* 21 -14])^(crc_i[15]&ahead[1023-32* 21 -15])^(crc_i[16]&ahead[1023-32* 21 -16])^(crc_i[17]&ahead[1023-32* 21 -17])^(crc_i[18]&ahead[1023-32* 21 -18])^(crc_i[19]&ahead[1023-32* 21 -19])^(crc_i[20]&ahead[1023-32* 21 -20])^(crc_i[21]&ahead[1023-32* 21 -21])^(crc_i[22]&ahead[1023-32* 21 -22])^(crc_i[23]&ahead[1023-32* 21 -23])^(crc_i[24]&ahead[1023-32* 21 -24])^(crc_i[25]&ahead[1023-32* 21 -25])^(crc_i[26]&ahead[1023-32* 21 -26])^(crc_i[27]&ahead[1023-32* 21 -27])^(crc_i[28]&ahead[1023-32* 21 -28])^(crc_i[29]&ahead[1023-32* 21 -29])^(crc_i[30]&ahead[1023-32* 21 -30])^(crc_i[31]&ahead[1023-32* 21 -31]);
// assign test[22] =    (crc_i[0]&ahead[1023-32* 22 ])^(crc_i[1]&ahead[1023-32* 22 -1])^(crc_i[2]&ahead[1023-32*22 -2 ])^(crc_i[3]&ahead[1023-32* 22 -3])^(crc_i[4]&ahead[1023-32* 22 -4])^(crc_i[5]&ahead[1023-32* 22 -5])^(crc_i[6]&ahead[1023-32* 22 -6])^(crc_i[7]&ahead[1023-32* 22 -7])^(crc_i[8]&ahead[1023-32* 22 -8])^(crc_i[9]&ahead[1023-32* 22 -9])^(crc_i[10]&ahead[1023-32* 22 -10])^(crc_i[11]&ahead[1023-32* 22 -11])^(crc_i[12]&ahead[1023-32* 22 -12])^(crc_i[13]&ahead[1023-32* 22 -13])^(crc_i[14]&ahead[1023-32* 22 -14])^(crc_i[15]&ahead[1023-32* 22 -15])^(crc_i[16]&ahead[1023-32* 22 -16])^(crc_i[17]&ahead[1023-32* 22 -17])^(crc_i[18]&ahead[1023-32* 22 -18])^(crc_i[19]&ahead[1023-32* 22 -19])^(crc_i[20]&ahead[1023-32* 22 -20])^(crc_i[21]&ahead[1023-32* 22 -21])^(crc_i[22]&ahead[1023-32* 22 -22])^(crc_i[23]&ahead[1023-32* 22 -23])^(crc_i[24]&ahead[1023-32* 22 -24])^(crc_i[25]&ahead[1023-32* 22 -25])^(crc_i[26]&ahead[1023-32* 22 -26])^(crc_i[27]&ahead[1023-32* 22 -27])^(crc_i[28]&ahead[1023-32* 22 -28])^(crc_i[29]&ahead[1023-32* 22 -29])^(crc_i[30]&ahead[1023-32* 22 -30])^(crc_i[31]&ahead[1023-32* 22 -31]);
// assign test[23] =    (crc_i[0]&ahead[1023-32* 23 ])^(crc_i[1]&ahead[1023-32* 23 -1])^(crc_i[2]&ahead[1023-32*23 -2 ])^(crc_i[3]&ahead[1023-32* 23 -3])^(crc_i[4]&ahead[1023-32* 23 -4])^(crc_i[5]&ahead[1023-32* 23 -5])^(crc_i[6]&ahead[1023-32* 23 -6])^(crc_i[7]&ahead[1023-32* 23 -7])^(crc_i[8]&ahead[1023-32* 23 -8])^(crc_i[9]&ahead[1023-32* 23 -9])^(crc_i[10]&ahead[1023-32* 23 -10])^(crc_i[11]&ahead[1023-32* 23 -11])^(crc_i[12]&ahead[1023-32* 23 -12])^(crc_i[13]&ahead[1023-32* 23 -13])^(crc_i[14]&ahead[1023-32* 23 -14])^(crc_i[15]&ahead[1023-32* 23 -15])^(crc_i[16]&ahead[1023-32* 23 -16])^(crc_i[17]&ahead[1023-32* 23 -17])^(crc_i[18]&ahead[1023-32* 23 -18])^(crc_i[19]&ahead[1023-32* 23 -19])^(crc_i[20]&ahead[1023-32* 23 -20])^(crc_i[21]&ahead[1023-32* 23 -21])^(crc_i[22]&ahead[1023-32* 23 -22])^(crc_i[23]&ahead[1023-32* 23 -23])^(crc_i[24]&ahead[1023-32* 23 -24])^(crc_i[25]&ahead[1023-32* 23 -25])^(crc_i[26]&ahead[1023-32* 23 -26])^(crc_i[27]&ahead[1023-32* 23 -27])^(crc_i[28]&ahead[1023-32* 23 -28])^(crc_i[29]&ahead[1023-32* 23 -29])^(crc_i[30]&ahead[1023-32* 23 -30])^(crc_i[31]&ahead[1023-32* 23 -31]);
// assign test[24] =    (crc_i[0]&ahead[1023-32* 24 ])^(crc_i[1]&ahead[1023-32* 24 -1])^(crc_i[2]&ahead[1023-32*24 -2 ])^(crc_i[3]&ahead[1023-32* 24 -3])^(crc_i[4]&ahead[1023-32* 24 -4])^(crc_i[5]&ahead[1023-32* 24 -5])^(crc_i[6]&ahead[1023-32* 24 -6])^(crc_i[7]&ahead[1023-32* 24 -7])^(crc_i[8]&ahead[1023-32* 24 -8])^(crc_i[9]&ahead[1023-32* 24 -9])^(crc_i[10]&ahead[1023-32* 24 -10])^(crc_i[11]&ahead[1023-32* 24 -11])^(crc_i[12]&ahead[1023-32* 24 -12])^(crc_i[13]&ahead[1023-32* 24 -13])^(crc_i[14]&ahead[1023-32* 24 -14])^(crc_i[15]&ahead[1023-32* 24 -15])^(crc_i[16]&ahead[1023-32* 24 -16])^(crc_i[17]&ahead[1023-32* 24 -17])^(crc_i[18]&ahead[1023-32* 24 -18])^(crc_i[19]&ahead[1023-32* 24 -19])^(crc_i[20]&ahead[1023-32* 24 -20])^(crc_i[21]&ahead[1023-32* 24 -21])^(crc_i[22]&ahead[1023-32* 24 -22])^(crc_i[23]&ahead[1023-32* 24 -23])^(crc_i[24]&ahead[1023-32* 24 -24])^(crc_i[25]&ahead[1023-32* 24 -25])^(crc_i[26]&ahead[1023-32* 24 -26])^(crc_i[27]&ahead[1023-32* 24 -27])^(crc_i[28]&ahead[1023-32* 24 -28])^(crc_i[29]&ahead[1023-32* 24 -29])^(crc_i[30]&ahead[1023-32* 24 -30])^(crc_i[31]&ahead[1023-32* 24 -31]);
// assign test[25] =    (crc_i[0]&ahead[1023-32* 25 ])^(crc_i[1]&ahead[1023-32* 25 -1])^(crc_i[2]&ahead[1023-32*25 -2 ])^(crc_i[3]&ahead[1023-32* 25 -3])^(crc_i[4]&ahead[1023-32* 25 -4])^(crc_i[5]&ahead[1023-32* 25 -5])^(crc_i[6]&ahead[1023-32* 25 -6])^(crc_i[7]&ahead[1023-32* 25 -7])^(crc_i[8]&ahead[1023-32* 25 -8])^(crc_i[9]&ahead[1023-32* 25 -9])^(crc_i[10]&ahead[1023-32* 25 -10])^(crc_i[11]&ahead[1023-32* 25 -11])^(crc_i[12]&ahead[1023-32* 25 -12])^(crc_i[13]&ahead[1023-32* 25 -13])^(crc_i[14]&ahead[1023-32* 25 -14])^(crc_i[15]&ahead[1023-32* 25 -15])^(crc_i[16]&ahead[1023-32* 25 -16])^(crc_i[17]&ahead[1023-32* 25 -17])^(crc_i[18]&ahead[1023-32* 25 -18])^(crc_i[19]&ahead[1023-32* 25 -19])^(crc_i[20]&ahead[1023-32* 25 -20])^(crc_i[21]&ahead[1023-32* 25 -21])^(crc_i[22]&ahead[1023-32* 25 -22])^(crc_i[23]&ahead[1023-32* 25 -23])^(crc_i[24]&ahead[1023-32* 25 -24])^(crc_i[25]&ahead[1023-32* 25 -25])^(crc_i[26]&ahead[1023-32* 25 -26])^(crc_i[27]&ahead[1023-32* 25 -27])^(crc_i[28]&ahead[1023-32* 25 -28])^(crc_i[29]&ahead[1023-32* 25 -29])^(crc_i[30]&ahead[1023-32* 25 -30])^(crc_i[31]&ahead[1023-32* 25 -31]);
// assign test[26] =    (crc_i[0]&ahead[1023-32* 26 ])^(crc_i[1]&ahead[1023-32* 26 -1])^(crc_i[2]&ahead[1023-32*26 -2 ])^(crc_i[3]&ahead[1023-32* 26 -3])^(crc_i[4]&ahead[1023-32* 26 -4])^(crc_i[5]&ahead[1023-32* 26 -5])^(crc_i[6]&ahead[1023-32* 26 -6])^(crc_i[7]&ahead[1023-32* 26 -7])^(crc_i[8]&ahead[1023-32* 26 -8])^(crc_i[9]&ahead[1023-32* 26 -9])^(crc_i[10]&ahead[1023-32* 26 -10])^(crc_i[11]&ahead[1023-32* 26 -11])^(crc_i[12]&ahead[1023-32* 26 -12])^(crc_i[13]&ahead[1023-32* 26 -13])^(crc_i[14]&ahead[1023-32* 26 -14])^(crc_i[15]&ahead[1023-32* 26 -15])^(crc_i[16]&ahead[1023-32* 26 -16])^(crc_i[17]&ahead[1023-32* 26 -17])^(crc_i[18]&ahead[1023-32* 26 -18])^(crc_i[19]&ahead[1023-32* 26 -19])^(crc_i[20]&ahead[1023-32* 26 -20])^(crc_i[21]&ahead[1023-32* 26 -21])^(crc_i[22]&ahead[1023-32* 26 -22])^(crc_i[23]&ahead[1023-32* 26 -23])^(crc_i[24]&ahead[1023-32* 26 -24])^(crc_i[25]&ahead[1023-32* 26 -25])^(crc_i[26]&ahead[1023-32* 26 -26])^(crc_i[27]&ahead[1023-32* 26 -27])^(crc_i[28]&ahead[1023-32* 26 -28])^(crc_i[29]&ahead[1023-32* 26 -29])^(crc_i[30]&ahead[1023-32* 26 -30])^(crc_i[31]&ahead[1023-32* 26 -31]);
// assign test[27] =    (crc_i[0]&ahead[1023-32* 27 ])^(crc_i[1]&ahead[1023-32* 27 -1])^(crc_i[2]&ahead[1023-32*27 -2 ])^(crc_i[3]&ahead[1023-32* 27 -3])^(crc_i[4]&ahead[1023-32* 27 -4])^(crc_i[5]&ahead[1023-32* 27 -5])^(crc_i[6]&ahead[1023-32* 27 -6])^(crc_i[7]&ahead[1023-32* 27 -7])^(crc_i[8]&ahead[1023-32* 27 -8])^(crc_i[9]&ahead[1023-32* 27 -9])^(crc_i[10]&ahead[1023-32* 27 -10])^(crc_i[11]&ahead[1023-32* 27 -11])^(crc_i[12]&ahead[1023-32* 27 -12])^(crc_i[13]&ahead[1023-32* 27 -13])^(crc_i[14]&ahead[1023-32* 27 -14])^(crc_i[15]&ahead[1023-32* 27 -15])^(crc_i[16]&ahead[1023-32* 27 -16])^(crc_i[17]&ahead[1023-32* 27 -17])^(crc_i[18]&ahead[1023-32* 27 -18])^(crc_i[19]&ahead[1023-32* 27 -19])^(crc_i[20]&ahead[1023-32* 27 -20])^(crc_i[21]&ahead[1023-32* 27 -21])^(crc_i[22]&ahead[1023-32* 27 -22])^(crc_i[23]&ahead[1023-32* 27 -23])^(crc_i[24]&ahead[1023-32* 27 -24])^(crc_i[25]&ahead[1023-32* 27 -25])^(crc_i[26]&ahead[1023-32* 27 -26])^(crc_i[27]&ahead[1023-32* 27 -27])^(crc_i[28]&ahead[1023-32* 27 -28])^(crc_i[29]&ahead[1023-32* 27 -29])^(crc_i[30]&ahead[1023-32* 27 -30])^(crc_i[31]&ahead[1023-32* 27 -31]);
// assign test[28] =    (crc_i[0]&ahead[1023-32* 28 ])^(crc_i[1]&ahead[1023-32* 28 -1])^(crc_i[2]&ahead[1023-32*28 -2 ])^(crc_i[3]&ahead[1023-32* 28 -3])^(crc_i[4]&ahead[1023-32* 28 -4])^(crc_i[5]&ahead[1023-32* 28 -5])^(crc_i[6]&ahead[1023-32* 28 -6])^(crc_i[7]&ahead[1023-32* 28 -7])^(crc_i[8]&ahead[1023-32* 28 -8])^(crc_i[9]&ahead[1023-32* 28 -9])^(crc_i[10]&ahead[1023-32* 28 -10])^(crc_i[11]&ahead[1023-32* 28 -11])^(crc_i[12]&ahead[1023-32* 28 -12])^(crc_i[13]&ahead[1023-32* 28 -13])^(crc_i[14]&ahead[1023-32* 28 -14])^(crc_i[15]&ahead[1023-32* 28 -15])^(crc_i[16]&ahead[1023-32* 28 -16])^(crc_i[17]&ahead[1023-32* 28 -17])^(crc_i[18]&ahead[1023-32* 28 -18])^(crc_i[19]&ahead[1023-32* 28 -19])^(crc_i[20]&ahead[1023-32* 28 -20])^(crc_i[21]&ahead[1023-32* 28 -21])^(crc_i[22]&ahead[1023-32* 28 -22])^(crc_i[23]&ahead[1023-32* 28 -23])^(crc_i[24]&ahead[1023-32* 28 -24])^(crc_i[25]&ahead[1023-32* 28 -25])^(crc_i[26]&ahead[1023-32* 28 -26])^(crc_i[27]&ahead[1023-32* 28 -27])^(crc_i[28]&ahead[1023-32* 28 -28])^(crc_i[29]&ahead[1023-32* 28 -29])^(crc_i[30]&ahead[1023-32* 28 -30])^(crc_i[31]&ahead[1023-32* 28 -31]);
// assign test[29] =    (crc_i[0]&ahead[1023-32* 29 ])^(crc_i[1]&ahead[1023-32* 29 -1])^(crc_i[2]&ahead[1023-32*29 -2 ])^(crc_i[3]&ahead[1023-32* 29 -3])^(crc_i[4]&ahead[1023-32* 29 -4])^(crc_i[5]&ahead[1023-32* 29 -5])^(crc_i[6]&ahead[1023-32* 29 -6])^(crc_i[7]&ahead[1023-32* 29 -7])^(crc_i[8]&ahead[1023-32* 29 -8])^(crc_i[9]&ahead[1023-32* 29 -9])^(crc_i[10]&ahead[1023-32* 29 -10])^(crc_i[11]&ahead[1023-32* 29 -11])^(crc_i[12]&ahead[1023-32* 29 -12])^(crc_i[13]&ahead[1023-32* 29 -13])^(crc_i[14]&ahead[1023-32* 29 -14])^(crc_i[15]&ahead[1023-32* 29 -15])^(crc_i[16]&ahead[1023-32* 29 -16])^(crc_i[17]&ahead[1023-32* 29 -17])^(crc_i[18]&ahead[1023-32* 29 -18])^(crc_i[19]&ahead[1023-32* 29 -19])^(crc_i[20]&ahead[1023-32* 29 -20])^(crc_i[21]&ahead[1023-32* 29 -21])^(crc_i[22]&ahead[1023-32* 29 -22])^(crc_i[23]&ahead[1023-32* 29 -23])^(crc_i[24]&ahead[1023-32* 29 -24])^(crc_i[25]&ahead[1023-32* 29 -25])^(crc_i[26]&ahead[1023-32* 29 -26])^(crc_i[27]&ahead[1023-32* 29 -27])^(crc_i[28]&ahead[1023-32* 29 -28])^(crc_i[29]&ahead[1023-32* 29 -29])^(crc_i[30]&ahead[1023-32* 29 -30])^(crc_i[31]&ahead[1023-32* 29 -31]);
// assign test[30] =    (crc_i[0]&ahead[1023-32* 30 ])^(crc_i[1]&ahead[1023-32* 30 -1])^(crc_i[2]&ahead[1023-32*30 -2 ])^(crc_i[3]&ahead[1023-32* 30 -3])^(crc_i[4]&ahead[1023-32* 30 -4])^(crc_i[5]&ahead[1023-32* 30 -5])^(crc_i[6]&ahead[1023-32* 30 -6])^(crc_i[7]&ahead[1023-32* 30 -7])^(crc_i[8]&ahead[1023-32* 30 -8])^(crc_i[9]&ahead[1023-32* 30 -9])^(crc_i[10]&ahead[1023-32* 30 -10])^(crc_i[11]&ahead[1023-32* 30 -11])^(crc_i[12]&ahead[1023-32* 30 -12])^(crc_i[13]&ahead[1023-32* 30 -13])^(crc_i[14]&ahead[1023-32* 30 -14])^(crc_i[15]&ahead[1023-32* 30 -15])^(crc_i[16]&ahead[1023-32* 30 -16])^(crc_i[17]&ahead[1023-32* 30 -17])^(crc_i[18]&ahead[1023-32* 30 -18])^(crc_i[19]&ahead[1023-32* 30 -19])^(crc_i[20]&ahead[1023-32* 30 -20])^(crc_i[21]&ahead[1023-32* 30 -21])^(crc_i[22]&ahead[1023-32* 30 -22])^(crc_i[23]&ahead[1023-32* 30 -23])^(crc_i[24]&ahead[1023-32* 30 -24])^(crc_i[25]&ahead[1023-32* 30 -25])^(crc_i[26]&ahead[1023-32* 30 -26])^(crc_i[27]&ahead[1023-32* 30 -27])^(crc_i[28]&ahead[1023-32* 30 -28])^(crc_i[29]&ahead[1023-32* 30 -29])^(crc_i[30]&ahead[1023-32* 30 -30])^(crc_i[31]&ahead[1023-32* 30 -31]);
// assign test[31] =    (crc_i[0]&ahead[1023-32* 31 ])^(crc_i[1]&ahead[1023-32* 31 -1])^(crc_i[2]&ahead[1023-32*31 -2 ])^(crc_i[3]&ahead[1023-32* 31 -3])^(crc_i[4]&ahead[1023-32* 31 -4])^(crc_i[5]&ahead[1023-32* 31 -5])^(crc_i[6]&ahead[1023-32* 31 -6])^(crc_i[7]&ahead[1023-32* 31 -7])^(crc_i[8]&ahead[1023-32* 31 -8])^(crc_i[9]&ahead[1023-32* 31 -9])^(crc_i[10]&ahead[1023-32* 31 -10])^(crc_i[11]&ahead[1023-32* 31 -11])^(crc_i[12]&ahead[1023-32* 31 -12])^(crc_i[13]&ahead[1023-32* 31 -13])^(crc_i[14]&ahead[1023-32* 31 -14])^(crc_i[15]&ahead[1023-32* 31 -15])^(crc_i[16]&ahead[1023-32* 31 -16])^(crc_i[17]&ahead[1023-32* 31 -17])^(crc_i[18]&ahead[1023-32* 31 -18])^(crc_i[19]&ahead[1023-32* 31 -19])^(crc_i[20]&ahead[1023-32* 31 -20])^(crc_i[21]&ahead[1023-32* 31 -21])^(crc_i[22]&ahead[1023-32* 31 -22])^(crc_i[23]&ahead[1023-32* 31 -23])^(crc_i[24]&ahead[1023-32* 31 -24])^(crc_i[25]&ahead[1023-32* 31 -25])^(crc_i[26]&ahead[1023-32* 31 -26])^(crc_i[27]&ahead[1023-32* 31 -27])^(crc_i[28]&ahead[1023-32* 31 -28])^(crc_i[29]&ahead[1023-32* 31 -29])^(crc_i[30]&ahead[1023-32* 31 -30])^(crc_i[31]&ahead[1023-32* 31 -31]);

// wire [31:0] test_wire ;


// assign test_wire[0 ] = (crc_i[0]&ahead[1023-32* 31 ]) ^(crc_i[1]&ahead[1023-32* 31 -1]) ^(crc_i[2]&ahead[1023-32* -2 ])^(crc_i[3]&ahead[1023-32* 31 -3])^(crc_i[4]&ahead[1023-32* 31 -4])^(crc_i[5]&ahead[1023-32* 31 -5])^(crc_i[6]&ahead[1023-32* 31 -6])^(crc_i[7]&ahead[1023-32* 31 -7])^(crc_i[8]&ahead[1023-32* 31 -8]) ; 
// assign test_wire[1 ] = (crc_i[0]&ahead[1023-32* 31 ]) ^(crc_i[1]&ahead[1023-32* 31 -1]) ^(crc_i[2]&ahead[1023-32* -2 ])^(crc_i[3]&ahead[1023-32* 31 -3])^(crc_i[4]&ahead[1023-32* 31 -4])^(crc_i[5]&ahead[1023-32* 31 -5])^(crc_i[6]&ahead[1023-32* 31 -6])^(crc_i[7]&ahead[1023-32* 31 -7]) ;
// assign test_wire[2 ] = (crc_i[0]&ahead[1023-32* 31 ]) ^(crc_i[1]&ahead[1023-32* 31 -1]) ^(crc_i[2]&ahead[1023-32* -2 ])^(crc_i[3]&ahead[1023-32* 31 -3])^(crc_i[4]&ahead[1023-32* 31 -4])^(crc_i[5]&ahead[1023-32* 31 -5])^(crc_i[6]&ahead[1023-32* 31 -6]) ;
// assign test_wire[3 ] = (crc_i[0]&ahead[1023-32* 31 ]) ^(crc_i[1]&ahead[1023-32* 31 -1]) ^(crc_i[2]&ahead[1023-32* -2 ])^(crc_i[3]&ahead[1023-32* 31 -3])^(crc_i[4]&ahead[1023-32* 31 -4])^(crc_i[5]&ahead[1023-32* 31 -5]) ;
// assign test_wire[4 ] = (crc_i[0]&ahead[1023-32* 31 ]) ^(crc_i[1]&ahead[1023-32* 31 -1]) ^(crc_i[2]&ahead[1023-32* -2 ])^(crc_i[3]&ahead[1023-32* 31 -3])^(crc_i[4]&ahead[1023-32* 31 -4]) ;
// assign test_wire[5 ] = (crc_i[0]&ahead[1023-32* 31 ]) ^(crc_i[1]&ahead[1023-32* 31 -1]) ^(crc_i[2]&ahead[1023-32* -2 ])^(crc_i[3]&ahead[1023-32* 31 -3]) ;
// assign test_wire[6 ] = (crc_i[0]&ahead[1023-32* 31 ]) ^(crc_i[1]&ahead[1023-32* 31 -1]) ^(crc_i[2]&ahead[1023-32* -2 ]) ;
// assign test_wire[7 ] = (crc_i[0]&ahead[1023-32* 31 ]) ^(crc_i[1]&ahead[1023-32* 31 -1]) ;
// assign test_wire[8 ] = (crc_i[0]&ahead[1023-32* 31 ]) ;



assign ahead[0 ] =    (crc_i[0]&AHEAD_POLY[1023-32* 0  ])^(crc_i[1]&AHEAD_POLY[1023-32* 0  -1])^(crc_i[2]&AHEAD_POLY[1023-32*0  -2 ])^(crc_i[3]&AHEAD_POLY[1023-32* 0  -3])^(crc_i[4]&AHEAD_POLY[1023-32* 0  -4])^(crc_i[5]&AHEAD_POLY[1023-32* 0  -5])^(crc_i[6]&AHEAD_POLY[1023-32* 0  -6])^(crc_i[7]&AHEAD_POLY[1023-32* 0  -7])^(crc_i[8]&AHEAD_POLY[1023-32* 0  -8])^(crc_i[9]&AHEAD_POLY[1023-32* 0  -9])^(crc_i[10]&AHEAD_POLY[1023-32* 0  -10])^(crc_i[11]&AHEAD_POLY[1023-32* 0  -11])^(crc_i[12]&AHEAD_POLY[1023-32* 0  -12])^(crc_i[13]&AHEAD_POLY[1023-32* 0  -13])^(crc_i[14]&AHEAD_POLY[1023-32* 0  -14])^(crc_i[15]&AHEAD_POLY[1023-32* 0  -15])^(crc_i[16]&AHEAD_POLY[1023-32* 0  -16])^(crc_i[17]&AHEAD_POLY[1023-32* 0  -17])^(crc_i[18]&AHEAD_POLY[1023-32* 0  -18])^(crc_i[19]&AHEAD_POLY[1023-32* 0  -19])^(crc_i[20]&AHEAD_POLY[1023-32* 0  -20])^(crc_i[21]&AHEAD_POLY[1023-32* 0  -21])^(crc_i[22]&AHEAD_POLY[1023-32* 0  -22])^(crc_i[23]&AHEAD_POLY[1023-32* 0  -23])^(crc_i[24]&AHEAD_POLY[1023-32* 0  -24])^(crc_i[25]&AHEAD_POLY[1023-32* 0  -25])^(crc_i[26]&AHEAD_POLY[1023-32* 0  -26])^(crc_i[27]&AHEAD_POLY[1023-32* 0  -27])^(crc_i[28]&AHEAD_POLY[1023-32* 0  -28])^(crc_i[29]&AHEAD_POLY[1023-32* 0  -29])^(crc_i[30]&AHEAD_POLY[1023-32* 0  -30])^(crc_i[31]&AHEAD_POLY[1023-32* 0  -31]);
assign ahead[1 ] =    (crc_i[0]&AHEAD_POLY[1023-32* 1  ])^(crc_i[1]&AHEAD_POLY[1023-32* 1  -1])^(crc_i[2]&AHEAD_POLY[1023-32*1  -2 ])^(crc_i[3]&AHEAD_POLY[1023-32* 1  -3])^(crc_i[4]&AHEAD_POLY[1023-32* 1  -4])^(crc_i[5]&AHEAD_POLY[1023-32* 1  -5])^(crc_i[6]&AHEAD_POLY[1023-32* 1  -6])^(crc_i[7]&AHEAD_POLY[1023-32* 1  -7])^(crc_i[8]&AHEAD_POLY[1023-32* 1  -8])^(crc_i[9]&AHEAD_POLY[1023-32* 1  -9])^(crc_i[10]&AHEAD_POLY[1023-32* 1  -10])^(crc_i[11]&AHEAD_POLY[1023-32* 1  -11])^(crc_i[12]&AHEAD_POLY[1023-32* 1  -12])^(crc_i[13]&AHEAD_POLY[1023-32* 1  -13])^(crc_i[14]&AHEAD_POLY[1023-32* 1  -14])^(crc_i[15]&AHEAD_POLY[1023-32* 1  -15])^(crc_i[16]&AHEAD_POLY[1023-32* 1  -16])^(crc_i[17]&AHEAD_POLY[1023-32* 1  -17])^(crc_i[18]&AHEAD_POLY[1023-32* 1  -18])^(crc_i[19]&AHEAD_POLY[1023-32* 1  -19])^(crc_i[20]&AHEAD_POLY[1023-32* 1  -20])^(crc_i[21]&AHEAD_POLY[1023-32* 1  -21])^(crc_i[22]&AHEAD_POLY[1023-32* 1  -22])^(crc_i[23]&AHEAD_POLY[1023-32* 1  -23])^(crc_i[24]&AHEAD_POLY[1023-32* 1  -24])^(crc_i[25]&AHEAD_POLY[1023-32* 1  -25])^(crc_i[26]&AHEAD_POLY[1023-32* 1  -26])^(crc_i[27]&AHEAD_POLY[1023-32* 1  -27])^(crc_i[28]&AHEAD_POLY[1023-32* 1  -28])^(crc_i[29]&AHEAD_POLY[1023-32* 1  -29])^(crc_i[30]&AHEAD_POLY[1023-32* 1  -30])^(crc_i[31]&AHEAD_POLY[1023-32* 1  -31]);
assign ahead[2 ] =    (crc_i[0]&AHEAD_POLY[1023-32* 2  ])^(crc_i[1]&AHEAD_POLY[1023-32* 2  -1])^(crc_i[2]&AHEAD_POLY[1023-32*2  -2 ])^(crc_i[3]&AHEAD_POLY[1023-32* 2  -3])^(crc_i[4]&AHEAD_POLY[1023-32* 2  -4])^(crc_i[5]&AHEAD_POLY[1023-32* 2  -5])^(crc_i[6]&AHEAD_POLY[1023-32* 2  -6])^(crc_i[7]&AHEAD_POLY[1023-32* 2  -7])^(crc_i[8]&AHEAD_POLY[1023-32* 2  -8])^(crc_i[9]&AHEAD_POLY[1023-32* 2  -9])^(crc_i[10]&AHEAD_POLY[1023-32* 2  -10])^(crc_i[11]&AHEAD_POLY[1023-32* 2  -11])^(crc_i[12]&AHEAD_POLY[1023-32* 2  -12])^(crc_i[13]&AHEAD_POLY[1023-32* 2  -13])^(crc_i[14]&AHEAD_POLY[1023-32* 2  -14])^(crc_i[15]&AHEAD_POLY[1023-32* 2  -15])^(crc_i[16]&AHEAD_POLY[1023-32* 2  -16])^(crc_i[17]&AHEAD_POLY[1023-32* 2  -17])^(crc_i[18]&AHEAD_POLY[1023-32* 2  -18])^(crc_i[19]&AHEAD_POLY[1023-32* 2  -19])^(crc_i[20]&AHEAD_POLY[1023-32* 2  -20])^(crc_i[21]&AHEAD_POLY[1023-32* 2  -21])^(crc_i[22]&AHEAD_POLY[1023-32* 2  -22])^(crc_i[23]&AHEAD_POLY[1023-32* 2  -23])^(crc_i[24]&AHEAD_POLY[1023-32* 2  -24])^(crc_i[25]&AHEAD_POLY[1023-32* 2  -25])^(crc_i[26]&AHEAD_POLY[1023-32* 2  -26])^(crc_i[27]&AHEAD_POLY[1023-32* 2  -27])^(crc_i[28]&AHEAD_POLY[1023-32* 2  -28])^(crc_i[29]&AHEAD_POLY[1023-32* 2  -29])^(crc_i[30]&AHEAD_POLY[1023-32* 2  -30])^(crc_i[31]&AHEAD_POLY[1023-32* 2  -31]);
assign ahead[3 ] =    (crc_i[0]&AHEAD_POLY[1023-32* 3  ])^(crc_i[1]&AHEAD_POLY[1023-32* 3  -1])^(crc_i[2]&AHEAD_POLY[1023-32*3  -2 ])^(crc_i[3]&AHEAD_POLY[1023-32* 3  -3])^(crc_i[4]&AHEAD_POLY[1023-32* 3  -4])^(crc_i[5]&AHEAD_POLY[1023-32* 3  -5])^(crc_i[6]&AHEAD_POLY[1023-32* 3  -6])^(crc_i[7]&AHEAD_POLY[1023-32* 3  -7])^(crc_i[8]&AHEAD_POLY[1023-32* 3  -8])^(crc_i[9]&AHEAD_POLY[1023-32* 3  -9])^(crc_i[10]&AHEAD_POLY[1023-32* 3  -10])^(crc_i[11]&AHEAD_POLY[1023-32* 3  -11])^(crc_i[12]&AHEAD_POLY[1023-32* 3  -12])^(crc_i[13]&AHEAD_POLY[1023-32* 3  -13])^(crc_i[14]&AHEAD_POLY[1023-32* 3  -14])^(crc_i[15]&AHEAD_POLY[1023-32* 3  -15])^(crc_i[16]&AHEAD_POLY[1023-32* 3  -16])^(crc_i[17]&AHEAD_POLY[1023-32* 3  -17])^(crc_i[18]&AHEAD_POLY[1023-32* 3  -18])^(crc_i[19]&AHEAD_POLY[1023-32* 3  -19])^(crc_i[20]&AHEAD_POLY[1023-32* 3  -20])^(crc_i[21]&AHEAD_POLY[1023-32* 3  -21])^(crc_i[22]&AHEAD_POLY[1023-32* 3  -22])^(crc_i[23]&AHEAD_POLY[1023-32* 3  -23])^(crc_i[24]&AHEAD_POLY[1023-32* 3  -24])^(crc_i[25]&AHEAD_POLY[1023-32* 3  -25])^(crc_i[26]&AHEAD_POLY[1023-32* 3  -26])^(crc_i[27]&AHEAD_POLY[1023-32* 3  -27])^(crc_i[28]&AHEAD_POLY[1023-32* 3  -28])^(crc_i[29]&AHEAD_POLY[1023-32* 3  -29])^(crc_i[30]&AHEAD_POLY[1023-32* 3  -30])^(crc_i[31]&AHEAD_POLY[1023-32* 3  -31]);
assign ahead[4 ] =    (crc_i[0]&AHEAD_POLY[1023-32* 4  ])^(crc_i[1]&AHEAD_POLY[1023-32* 4  -1])^(crc_i[2]&AHEAD_POLY[1023-32*4  -2 ])^(crc_i[3]&AHEAD_POLY[1023-32* 4  -3])^(crc_i[4]&AHEAD_POLY[1023-32* 4  -4])^(crc_i[5]&AHEAD_POLY[1023-32* 4  -5])^(crc_i[6]&AHEAD_POLY[1023-32* 4  -6])^(crc_i[7]&AHEAD_POLY[1023-32* 4  -7])^(crc_i[8]&AHEAD_POLY[1023-32* 4  -8])^(crc_i[9]&AHEAD_POLY[1023-32* 4  -9])^(crc_i[10]&AHEAD_POLY[1023-32* 4  -10])^(crc_i[11]&AHEAD_POLY[1023-32* 4  -11])^(crc_i[12]&AHEAD_POLY[1023-32* 4  -12])^(crc_i[13]&AHEAD_POLY[1023-32* 4  -13])^(crc_i[14]&AHEAD_POLY[1023-32* 4  -14])^(crc_i[15]&AHEAD_POLY[1023-32* 4  -15])^(crc_i[16]&AHEAD_POLY[1023-32* 4  -16])^(crc_i[17]&AHEAD_POLY[1023-32* 4  -17])^(crc_i[18]&AHEAD_POLY[1023-32* 4  -18])^(crc_i[19]&AHEAD_POLY[1023-32* 4  -19])^(crc_i[20]&AHEAD_POLY[1023-32* 4  -20])^(crc_i[21]&AHEAD_POLY[1023-32* 4  -21])^(crc_i[22]&AHEAD_POLY[1023-32* 4  -22])^(crc_i[23]&AHEAD_POLY[1023-32* 4  -23])^(crc_i[24]&AHEAD_POLY[1023-32* 4  -24])^(crc_i[25]&AHEAD_POLY[1023-32* 4  -25])^(crc_i[26]&AHEAD_POLY[1023-32* 4  -26])^(crc_i[27]&AHEAD_POLY[1023-32* 4  -27])^(crc_i[28]&AHEAD_POLY[1023-32* 4  -28])^(crc_i[29]&AHEAD_POLY[1023-32* 4  -29])^(crc_i[30]&AHEAD_POLY[1023-32* 4  -30])^(crc_i[31]&AHEAD_POLY[1023-32* 4  -31]);
assign ahead[5 ] =    (crc_i[0]&AHEAD_POLY[1023-32* 5  ])^(crc_i[1]&AHEAD_POLY[1023-32* 5  -1])^(crc_i[2]&AHEAD_POLY[1023-32*5  -2 ])^(crc_i[3]&AHEAD_POLY[1023-32* 5  -3])^(crc_i[4]&AHEAD_POLY[1023-32* 5  -4])^(crc_i[5]&AHEAD_POLY[1023-32* 5  -5])^(crc_i[6]&AHEAD_POLY[1023-32* 5  -6])^(crc_i[7]&AHEAD_POLY[1023-32* 5  -7])^(crc_i[8]&AHEAD_POLY[1023-32* 5  -8])^(crc_i[9]&AHEAD_POLY[1023-32* 5  -9])^(crc_i[10]&AHEAD_POLY[1023-32* 5  -10])^(crc_i[11]&AHEAD_POLY[1023-32* 5  -11])^(crc_i[12]&AHEAD_POLY[1023-32* 5  -12])^(crc_i[13]&AHEAD_POLY[1023-32* 5  -13])^(crc_i[14]&AHEAD_POLY[1023-32* 5  -14])^(crc_i[15]&AHEAD_POLY[1023-32* 5  -15])^(crc_i[16]&AHEAD_POLY[1023-32* 5  -16])^(crc_i[17]&AHEAD_POLY[1023-32* 5  -17])^(crc_i[18]&AHEAD_POLY[1023-32* 5  -18])^(crc_i[19]&AHEAD_POLY[1023-32* 5  -19])^(crc_i[20]&AHEAD_POLY[1023-32* 5  -20])^(crc_i[21]&AHEAD_POLY[1023-32* 5  -21])^(crc_i[22]&AHEAD_POLY[1023-32* 5  -22])^(crc_i[23]&AHEAD_POLY[1023-32* 5  -23])^(crc_i[24]&AHEAD_POLY[1023-32* 5  -24])^(crc_i[25]&AHEAD_POLY[1023-32* 5  -25])^(crc_i[26]&AHEAD_POLY[1023-32* 5  -26])^(crc_i[27]&AHEAD_POLY[1023-32* 5  -27])^(crc_i[28]&AHEAD_POLY[1023-32* 5  -28])^(crc_i[29]&AHEAD_POLY[1023-32* 5  -29])^(crc_i[30]&AHEAD_POLY[1023-32* 5  -30])^(crc_i[31]&AHEAD_POLY[1023-32* 5  -31]);
assign ahead[6 ] =    (crc_i[0]&AHEAD_POLY[1023-32* 6  ])^(crc_i[1]&AHEAD_POLY[1023-32* 6  -1])^(crc_i[2]&AHEAD_POLY[1023-32*6  -2 ])^(crc_i[3]&AHEAD_POLY[1023-32* 6  -3])^(crc_i[4]&AHEAD_POLY[1023-32* 6  -4])^(crc_i[5]&AHEAD_POLY[1023-32* 6  -5])^(crc_i[6]&AHEAD_POLY[1023-32* 6  -6])^(crc_i[7]&AHEAD_POLY[1023-32* 6  -7])^(crc_i[8]&AHEAD_POLY[1023-32* 6  -8])^(crc_i[9]&AHEAD_POLY[1023-32* 6  -9])^(crc_i[10]&AHEAD_POLY[1023-32* 6  -10])^(crc_i[11]&AHEAD_POLY[1023-32* 6  -11])^(crc_i[12]&AHEAD_POLY[1023-32* 6  -12])^(crc_i[13]&AHEAD_POLY[1023-32* 6  -13])^(crc_i[14]&AHEAD_POLY[1023-32* 6  -14])^(crc_i[15]&AHEAD_POLY[1023-32* 6  -15])^(crc_i[16]&AHEAD_POLY[1023-32* 6  -16])^(crc_i[17]&AHEAD_POLY[1023-32* 6  -17])^(crc_i[18]&AHEAD_POLY[1023-32* 6  -18])^(crc_i[19]&AHEAD_POLY[1023-32* 6  -19])^(crc_i[20]&AHEAD_POLY[1023-32* 6  -20])^(crc_i[21]&AHEAD_POLY[1023-32* 6  -21])^(crc_i[22]&AHEAD_POLY[1023-32* 6  -22])^(crc_i[23]&AHEAD_POLY[1023-32* 6  -23])^(crc_i[24]&AHEAD_POLY[1023-32* 6  -24])^(crc_i[25]&AHEAD_POLY[1023-32* 6  -25])^(crc_i[26]&AHEAD_POLY[1023-32* 6  -26])^(crc_i[27]&AHEAD_POLY[1023-32* 6  -27])^(crc_i[28]&AHEAD_POLY[1023-32* 6  -28])^(crc_i[29]&AHEAD_POLY[1023-32* 6  -29])^(crc_i[30]&AHEAD_POLY[1023-32* 6  -30])^(crc_i[31]&AHEAD_POLY[1023-32* 6  -31]);
assign ahead[7 ] =    (crc_i[0]&AHEAD_POLY[1023-32* 7  ])^(crc_i[1]&AHEAD_POLY[1023-32* 7  -1])^(crc_i[2]&AHEAD_POLY[1023-32*7  -2 ])^(crc_i[3]&AHEAD_POLY[1023-32* 7  -3])^(crc_i[4]&AHEAD_POLY[1023-32* 7  -4])^(crc_i[5]&AHEAD_POLY[1023-32* 7  -5])^(crc_i[6]&AHEAD_POLY[1023-32* 7  -6])^(crc_i[7]&AHEAD_POLY[1023-32* 7  -7])^(crc_i[8]&AHEAD_POLY[1023-32* 7  -8])^(crc_i[9]&AHEAD_POLY[1023-32* 7  -9])^(crc_i[10]&AHEAD_POLY[1023-32* 7  -10])^(crc_i[11]&AHEAD_POLY[1023-32* 7  -11])^(crc_i[12]&AHEAD_POLY[1023-32* 7  -12])^(crc_i[13]&AHEAD_POLY[1023-32* 7  -13])^(crc_i[14]&AHEAD_POLY[1023-32* 7  -14])^(crc_i[15]&AHEAD_POLY[1023-32* 7  -15])^(crc_i[16]&AHEAD_POLY[1023-32* 7  -16])^(crc_i[17]&AHEAD_POLY[1023-32* 7  -17])^(crc_i[18]&AHEAD_POLY[1023-32* 7  -18])^(crc_i[19]&AHEAD_POLY[1023-32* 7  -19])^(crc_i[20]&AHEAD_POLY[1023-32* 7  -20])^(crc_i[21]&AHEAD_POLY[1023-32* 7  -21])^(crc_i[22]&AHEAD_POLY[1023-32* 7  -22])^(crc_i[23]&AHEAD_POLY[1023-32* 7  -23])^(crc_i[24]&AHEAD_POLY[1023-32* 7  -24])^(crc_i[25]&AHEAD_POLY[1023-32* 7  -25])^(crc_i[26]&AHEAD_POLY[1023-32* 7  -26])^(crc_i[27]&AHEAD_POLY[1023-32* 7  -27])^(crc_i[28]&AHEAD_POLY[1023-32* 7  -28])^(crc_i[29]&AHEAD_POLY[1023-32* 7  -29])^(crc_i[30]&AHEAD_POLY[1023-32* 7  -30])^(crc_i[31]&AHEAD_POLY[1023-32* 7  -31]);
assign ahead[8 ] =    (crc_i[0]&AHEAD_POLY[1023-32* 8  ])^(crc_i[1]&AHEAD_POLY[1023-32* 8  -1])^(crc_i[2]&AHEAD_POLY[1023-32*8  -2 ])^(crc_i[3]&AHEAD_POLY[1023-32* 8  -3])^(crc_i[4]&AHEAD_POLY[1023-32* 8  -4])^(crc_i[5]&AHEAD_POLY[1023-32* 8  -5])^(crc_i[6]&AHEAD_POLY[1023-32* 8  -6])^(crc_i[7]&AHEAD_POLY[1023-32* 8  -7])^(crc_i[8]&AHEAD_POLY[1023-32* 8  -8])^(crc_i[9]&AHEAD_POLY[1023-32* 8  -9])^(crc_i[10]&AHEAD_POLY[1023-32* 8  -10])^(crc_i[11]&AHEAD_POLY[1023-32* 8  -11])^(crc_i[12]&AHEAD_POLY[1023-32* 8  -12])^(crc_i[13]&AHEAD_POLY[1023-32* 8  -13])^(crc_i[14]&AHEAD_POLY[1023-32* 8  -14])^(crc_i[15]&AHEAD_POLY[1023-32* 8  -15])^(crc_i[16]&AHEAD_POLY[1023-32* 8  -16])^(crc_i[17]&AHEAD_POLY[1023-32* 8  -17])^(crc_i[18]&AHEAD_POLY[1023-32* 8  -18])^(crc_i[19]&AHEAD_POLY[1023-32* 8  -19])^(crc_i[20]&AHEAD_POLY[1023-32* 8  -20])^(crc_i[21]&AHEAD_POLY[1023-32* 8  -21])^(crc_i[22]&AHEAD_POLY[1023-32* 8  -22])^(crc_i[23]&AHEAD_POLY[1023-32* 8  -23])^(crc_i[24]&AHEAD_POLY[1023-32* 8  -24])^(crc_i[25]&AHEAD_POLY[1023-32* 8  -25])^(crc_i[26]&AHEAD_POLY[1023-32* 8  -26])^(crc_i[27]&AHEAD_POLY[1023-32* 8  -27])^(crc_i[28]&AHEAD_POLY[1023-32* 8  -28])^(crc_i[29]&AHEAD_POLY[1023-32* 8  -29])^(crc_i[30]&AHEAD_POLY[1023-32* 8  -30])^(crc_i[31]&AHEAD_POLY[1023-32* 8  -31]);
assign ahead[9 ] =    (crc_i[0]&AHEAD_POLY[1023-32* 9  ])^(crc_i[1]&AHEAD_POLY[1023-32* 9  -1])^(crc_i[2]&AHEAD_POLY[1023-32*9  -2 ])^(crc_i[3]&AHEAD_POLY[1023-32* 9  -3])^(crc_i[4]&AHEAD_POLY[1023-32* 9  -4])^(crc_i[5]&AHEAD_POLY[1023-32* 9  -5])^(crc_i[6]&AHEAD_POLY[1023-32* 9  -6])^(crc_i[7]&AHEAD_POLY[1023-32* 9  -7])^(crc_i[8]&AHEAD_POLY[1023-32* 9  -8])^(crc_i[9]&AHEAD_POLY[1023-32* 9  -9])^(crc_i[10]&AHEAD_POLY[1023-32* 9  -10])^(crc_i[11]&AHEAD_POLY[1023-32* 9  -11])^(crc_i[12]&AHEAD_POLY[1023-32* 9  -12])^(crc_i[13]&AHEAD_POLY[1023-32* 9  -13])^(crc_i[14]&AHEAD_POLY[1023-32* 9  -14])^(crc_i[15]&AHEAD_POLY[1023-32* 9  -15])^(crc_i[16]&AHEAD_POLY[1023-32* 9  -16])^(crc_i[17]&AHEAD_POLY[1023-32* 9  -17])^(crc_i[18]&AHEAD_POLY[1023-32* 9  -18])^(crc_i[19]&AHEAD_POLY[1023-32* 9  -19])^(crc_i[20]&AHEAD_POLY[1023-32* 9  -20])^(crc_i[21]&AHEAD_POLY[1023-32* 9  -21])^(crc_i[22]&AHEAD_POLY[1023-32* 9  -22])^(crc_i[23]&AHEAD_POLY[1023-32* 9  -23])^(crc_i[24]&AHEAD_POLY[1023-32* 9  -24])^(crc_i[25]&AHEAD_POLY[1023-32* 9  -25])^(crc_i[26]&AHEAD_POLY[1023-32* 9  -26])^(crc_i[27]&AHEAD_POLY[1023-32* 9  -27])^(crc_i[28]&AHEAD_POLY[1023-32* 9  -28])^(crc_i[29]&AHEAD_POLY[1023-32* 9  -29])^(crc_i[30]&AHEAD_POLY[1023-32* 9  -30])^(crc_i[31]&AHEAD_POLY[1023-32* 9  -31]);
assign ahead[10] =    (crc_i[0]&AHEAD_POLY[1023-32* 10 ])^(crc_i[1]&AHEAD_POLY[1023-32* 10 -1])^(crc_i[2]&AHEAD_POLY[1023-32*10 -2 ])^(crc_i[3]&AHEAD_POLY[1023-32* 10 -3])^(crc_i[4]&AHEAD_POLY[1023-32* 10 -4])^(crc_i[5]&AHEAD_POLY[1023-32* 10 -5])^(crc_i[6]&AHEAD_POLY[1023-32* 10 -6])^(crc_i[7]&AHEAD_POLY[1023-32* 10 -7])^(crc_i[8]&AHEAD_POLY[1023-32* 10 -8])^(crc_i[9]&AHEAD_POLY[1023-32* 10 -9])^(crc_i[10]&AHEAD_POLY[1023-32* 10 -10])^(crc_i[11]&AHEAD_POLY[1023-32* 10 -11])^(crc_i[12]&AHEAD_POLY[1023-32* 10 -12])^(crc_i[13]&AHEAD_POLY[1023-32* 10 -13])^(crc_i[14]&AHEAD_POLY[1023-32* 10 -14])^(crc_i[15]&AHEAD_POLY[1023-32* 10 -15])^(crc_i[16]&AHEAD_POLY[1023-32* 10 -16])^(crc_i[17]&AHEAD_POLY[1023-32* 10 -17])^(crc_i[18]&AHEAD_POLY[1023-32* 10 -18])^(crc_i[19]&AHEAD_POLY[1023-32* 10 -19])^(crc_i[20]&AHEAD_POLY[1023-32* 10 -20])^(crc_i[21]&AHEAD_POLY[1023-32* 10 -21])^(crc_i[22]&AHEAD_POLY[1023-32* 10 -22])^(crc_i[23]&AHEAD_POLY[1023-32* 10 -23])^(crc_i[24]&AHEAD_POLY[1023-32* 10 -24])^(crc_i[25]&AHEAD_POLY[1023-32* 10 -25])^(crc_i[26]&AHEAD_POLY[1023-32* 10 -26])^(crc_i[27]&AHEAD_POLY[1023-32* 10 -27])^(crc_i[28]&AHEAD_POLY[1023-32* 10 -28])^(crc_i[29]&AHEAD_POLY[1023-32* 10 -29])^(crc_i[30]&AHEAD_POLY[1023-32* 10 -30])^(crc_i[31]&AHEAD_POLY[1023-32* 10 -31]);
assign ahead[11] =    (crc_i[0]&AHEAD_POLY[1023-32* 11 ])^(crc_i[1]&AHEAD_POLY[1023-32* 11 -1])^(crc_i[2]&AHEAD_POLY[1023-32*11 -2 ])^(crc_i[3]&AHEAD_POLY[1023-32* 11 -3])^(crc_i[4]&AHEAD_POLY[1023-32* 11 -4])^(crc_i[5]&AHEAD_POLY[1023-32* 11 -5])^(crc_i[6]&AHEAD_POLY[1023-32* 11 -6])^(crc_i[7]&AHEAD_POLY[1023-32* 11 -7])^(crc_i[8]&AHEAD_POLY[1023-32* 11 -8])^(crc_i[9]&AHEAD_POLY[1023-32* 11 -9])^(crc_i[10]&AHEAD_POLY[1023-32* 11 -10])^(crc_i[11]&AHEAD_POLY[1023-32* 11 -11])^(crc_i[12]&AHEAD_POLY[1023-32* 11 -12])^(crc_i[13]&AHEAD_POLY[1023-32* 11 -13])^(crc_i[14]&AHEAD_POLY[1023-32* 11 -14])^(crc_i[15]&AHEAD_POLY[1023-32* 11 -15])^(crc_i[16]&AHEAD_POLY[1023-32* 11 -16])^(crc_i[17]&AHEAD_POLY[1023-32* 11 -17])^(crc_i[18]&AHEAD_POLY[1023-32* 11 -18])^(crc_i[19]&AHEAD_POLY[1023-32* 11 -19])^(crc_i[20]&AHEAD_POLY[1023-32* 11 -20])^(crc_i[21]&AHEAD_POLY[1023-32* 11 -21])^(crc_i[22]&AHEAD_POLY[1023-32* 11 -22])^(crc_i[23]&AHEAD_POLY[1023-32* 11 -23])^(crc_i[24]&AHEAD_POLY[1023-32* 11 -24])^(crc_i[25]&AHEAD_POLY[1023-32* 11 -25])^(crc_i[26]&AHEAD_POLY[1023-32* 11 -26])^(crc_i[27]&AHEAD_POLY[1023-32* 11 -27])^(crc_i[28]&AHEAD_POLY[1023-32* 11 -28])^(crc_i[29]&AHEAD_POLY[1023-32* 11 -29])^(crc_i[30]&AHEAD_POLY[1023-32* 11 -30])^(crc_i[31]&AHEAD_POLY[1023-32* 11 -31]);
assign ahead[12] =    (crc_i[0]&AHEAD_POLY[1023-32* 12 ])^(crc_i[1]&AHEAD_POLY[1023-32* 12 -1])^(crc_i[2]&AHEAD_POLY[1023-32*12 -2 ])^(crc_i[3]&AHEAD_POLY[1023-32* 12 -3])^(crc_i[4]&AHEAD_POLY[1023-32* 12 -4])^(crc_i[5]&AHEAD_POLY[1023-32* 12 -5])^(crc_i[6]&AHEAD_POLY[1023-32* 12 -6])^(crc_i[7]&AHEAD_POLY[1023-32* 12 -7])^(crc_i[8]&AHEAD_POLY[1023-32* 12 -8])^(crc_i[9]&AHEAD_POLY[1023-32* 12 -9])^(crc_i[10]&AHEAD_POLY[1023-32* 12 -10])^(crc_i[11]&AHEAD_POLY[1023-32* 12 -11])^(crc_i[12]&AHEAD_POLY[1023-32* 12 -12])^(crc_i[13]&AHEAD_POLY[1023-32* 12 -13])^(crc_i[14]&AHEAD_POLY[1023-32* 12 -14])^(crc_i[15]&AHEAD_POLY[1023-32* 12 -15])^(crc_i[16]&AHEAD_POLY[1023-32* 12 -16])^(crc_i[17]&AHEAD_POLY[1023-32* 12 -17])^(crc_i[18]&AHEAD_POLY[1023-32* 12 -18])^(crc_i[19]&AHEAD_POLY[1023-32* 12 -19])^(crc_i[20]&AHEAD_POLY[1023-32* 12 -20])^(crc_i[21]&AHEAD_POLY[1023-32* 12 -21])^(crc_i[22]&AHEAD_POLY[1023-32* 12 -22])^(crc_i[23]&AHEAD_POLY[1023-32* 12 -23])^(crc_i[24]&AHEAD_POLY[1023-32* 12 -24])^(crc_i[25]&AHEAD_POLY[1023-32* 12 -25])^(crc_i[26]&AHEAD_POLY[1023-32* 12 -26])^(crc_i[27]&AHEAD_POLY[1023-32* 12 -27])^(crc_i[28]&AHEAD_POLY[1023-32* 12 -28])^(crc_i[29]&AHEAD_POLY[1023-32* 12 -29])^(crc_i[30]&AHEAD_POLY[1023-32* 12 -30])^(crc_i[31]&AHEAD_POLY[1023-32* 12 -31]);
assign ahead[13] =    (crc_i[0]&AHEAD_POLY[1023-32* 13 ])^(crc_i[1]&AHEAD_POLY[1023-32* 13 -1])^(crc_i[2]&AHEAD_POLY[1023-32*13 -2 ])^(crc_i[3]&AHEAD_POLY[1023-32* 13 -3])^(crc_i[4]&AHEAD_POLY[1023-32* 13 -4])^(crc_i[5]&AHEAD_POLY[1023-32* 13 -5])^(crc_i[6]&AHEAD_POLY[1023-32* 13 -6])^(crc_i[7]&AHEAD_POLY[1023-32* 13 -7])^(crc_i[8]&AHEAD_POLY[1023-32* 13 -8])^(crc_i[9]&AHEAD_POLY[1023-32* 13 -9])^(crc_i[10]&AHEAD_POLY[1023-32* 13 -10])^(crc_i[11]&AHEAD_POLY[1023-32* 13 -11])^(crc_i[12]&AHEAD_POLY[1023-32* 13 -12])^(crc_i[13]&AHEAD_POLY[1023-32* 13 -13])^(crc_i[14]&AHEAD_POLY[1023-32* 13 -14])^(crc_i[15]&AHEAD_POLY[1023-32* 13 -15])^(crc_i[16]&AHEAD_POLY[1023-32* 13 -16])^(crc_i[17]&AHEAD_POLY[1023-32* 13 -17])^(crc_i[18]&AHEAD_POLY[1023-32* 13 -18])^(crc_i[19]&AHEAD_POLY[1023-32* 13 -19])^(crc_i[20]&AHEAD_POLY[1023-32* 13 -20])^(crc_i[21]&AHEAD_POLY[1023-32* 13 -21])^(crc_i[22]&AHEAD_POLY[1023-32* 13 -22])^(crc_i[23]&AHEAD_POLY[1023-32* 13 -23])^(crc_i[24]&AHEAD_POLY[1023-32* 13 -24])^(crc_i[25]&AHEAD_POLY[1023-32* 13 -25])^(crc_i[26]&AHEAD_POLY[1023-32* 13 -26])^(crc_i[27]&AHEAD_POLY[1023-32* 13 -27])^(crc_i[28]&AHEAD_POLY[1023-32* 13 -28])^(crc_i[29]&AHEAD_POLY[1023-32* 13 -29])^(crc_i[30]&AHEAD_POLY[1023-32* 13 -30])^(crc_i[31]&AHEAD_POLY[1023-32* 13 -31]);
assign ahead[14] =    (crc_i[0]&AHEAD_POLY[1023-32* 14 ])^(crc_i[1]&AHEAD_POLY[1023-32* 14 -1])^(crc_i[2]&AHEAD_POLY[1023-32*14 -2 ])^(crc_i[3]&AHEAD_POLY[1023-32* 14 -3])^(crc_i[4]&AHEAD_POLY[1023-32* 14 -4])^(crc_i[5]&AHEAD_POLY[1023-32* 14 -5])^(crc_i[6]&AHEAD_POLY[1023-32* 14 -6])^(crc_i[7]&AHEAD_POLY[1023-32* 14 -7])^(crc_i[8]&AHEAD_POLY[1023-32* 14 -8])^(crc_i[9]&AHEAD_POLY[1023-32* 14 -9])^(crc_i[10]&AHEAD_POLY[1023-32* 14 -10])^(crc_i[11]&AHEAD_POLY[1023-32* 14 -11])^(crc_i[12]&AHEAD_POLY[1023-32* 14 -12])^(crc_i[13]&AHEAD_POLY[1023-32* 14 -13])^(crc_i[14]&AHEAD_POLY[1023-32* 14 -14])^(crc_i[15]&AHEAD_POLY[1023-32* 14 -15])^(crc_i[16]&AHEAD_POLY[1023-32* 14 -16])^(crc_i[17]&AHEAD_POLY[1023-32* 14 -17])^(crc_i[18]&AHEAD_POLY[1023-32* 14 -18])^(crc_i[19]&AHEAD_POLY[1023-32* 14 -19])^(crc_i[20]&AHEAD_POLY[1023-32* 14 -20])^(crc_i[21]&AHEAD_POLY[1023-32* 14 -21])^(crc_i[22]&AHEAD_POLY[1023-32* 14 -22])^(crc_i[23]&AHEAD_POLY[1023-32* 14 -23])^(crc_i[24]&AHEAD_POLY[1023-32* 14 -24])^(crc_i[25]&AHEAD_POLY[1023-32* 14 -25])^(crc_i[26]&AHEAD_POLY[1023-32* 14 -26])^(crc_i[27]&AHEAD_POLY[1023-32* 14 -27])^(crc_i[28]&AHEAD_POLY[1023-32* 14 -28])^(crc_i[29]&AHEAD_POLY[1023-32* 14 -29])^(crc_i[30]&AHEAD_POLY[1023-32* 14 -30])^(crc_i[31]&AHEAD_POLY[1023-32* 14 -31]);
assign ahead[15] =    (crc_i[0]&AHEAD_POLY[1023-32* 15 ])^(crc_i[1]&AHEAD_POLY[1023-32* 15 -1])^(crc_i[2]&AHEAD_POLY[1023-32*15 -2 ])^(crc_i[3]&AHEAD_POLY[1023-32* 15 -3])^(crc_i[4]&AHEAD_POLY[1023-32* 15 -4])^(crc_i[5]&AHEAD_POLY[1023-32* 15 -5])^(crc_i[6]&AHEAD_POLY[1023-32* 15 -6])^(crc_i[7]&AHEAD_POLY[1023-32* 15 -7])^(crc_i[8]&AHEAD_POLY[1023-32* 15 -8])^(crc_i[9]&AHEAD_POLY[1023-32* 15 -9])^(crc_i[10]&AHEAD_POLY[1023-32* 15 -10])^(crc_i[11]&AHEAD_POLY[1023-32* 15 -11])^(crc_i[12]&AHEAD_POLY[1023-32* 15 -12])^(crc_i[13]&AHEAD_POLY[1023-32* 15 -13])^(crc_i[14]&AHEAD_POLY[1023-32* 15 -14])^(crc_i[15]&AHEAD_POLY[1023-32* 15 -15])^(crc_i[16]&AHEAD_POLY[1023-32* 15 -16])^(crc_i[17]&AHEAD_POLY[1023-32* 15 -17])^(crc_i[18]&AHEAD_POLY[1023-32* 15 -18])^(crc_i[19]&AHEAD_POLY[1023-32* 15 -19])^(crc_i[20]&AHEAD_POLY[1023-32* 15 -20])^(crc_i[21]&AHEAD_POLY[1023-32* 15 -21])^(crc_i[22]&AHEAD_POLY[1023-32* 15 -22])^(crc_i[23]&AHEAD_POLY[1023-32* 15 -23])^(crc_i[24]&AHEAD_POLY[1023-32* 15 -24])^(crc_i[25]&AHEAD_POLY[1023-32* 15 -25])^(crc_i[26]&AHEAD_POLY[1023-32* 15 -26])^(crc_i[27]&AHEAD_POLY[1023-32* 15 -27])^(crc_i[28]&AHEAD_POLY[1023-32* 15 -28])^(crc_i[29]&AHEAD_POLY[1023-32* 15 -29])^(crc_i[30]&AHEAD_POLY[1023-32* 15 -30])^(crc_i[31]&AHEAD_POLY[1023-32* 15 -31]);
assign ahead[16] =    (crc_i[0]&AHEAD_POLY[1023-32* 16 ])^(crc_i[1]&AHEAD_POLY[1023-32* 16 -1])^(crc_i[2]&AHEAD_POLY[1023-32*16 -2 ])^(crc_i[3]&AHEAD_POLY[1023-32* 16 -3])^(crc_i[4]&AHEAD_POLY[1023-32* 16 -4])^(crc_i[5]&AHEAD_POLY[1023-32* 16 -5])^(crc_i[6]&AHEAD_POLY[1023-32* 16 -6])^(crc_i[7]&AHEAD_POLY[1023-32* 16 -7])^(crc_i[8]&AHEAD_POLY[1023-32* 16 -8])^(crc_i[9]&AHEAD_POLY[1023-32* 16 -9])^(crc_i[10]&AHEAD_POLY[1023-32* 16 -10])^(crc_i[11]&AHEAD_POLY[1023-32* 16 -11])^(crc_i[12]&AHEAD_POLY[1023-32* 16 -12])^(crc_i[13]&AHEAD_POLY[1023-32* 16 -13])^(crc_i[14]&AHEAD_POLY[1023-32* 16 -14])^(crc_i[15]&AHEAD_POLY[1023-32* 16 -15])^(crc_i[16]&AHEAD_POLY[1023-32* 16 -16])^(crc_i[17]&AHEAD_POLY[1023-32* 16 -17])^(crc_i[18]&AHEAD_POLY[1023-32* 16 -18])^(crc_i[19]&AHEAD_POLY[1023-32* 16 -19])^(crc_i[20]&AHEAD_POLY[1023-32* 16 -20])^(crc_i[21]&AHEAD_POLY[1023-32* 16 -21])^(crc_i[22]&AHEAD_POLY[1023-32* 16 -22])^(crc_i[23]&AHEAD_POLY[1023-32* 16 -23])^(crc_i[24]&AHEAD_POLY[1023-32* 16 -24])^(crc_i[25]&AHEAD_POLY[1023-32* 16 -25])^(crc_i[26]&AHEAD_POLY[1023-32* 16 -26])^(crc_i[27]&AHEAD_POLY[1023-32* 16 -27])^(crc_i[28]&AHEAD_POLY[1023-32* 16 -28])^(crc_i[29]&AHEAD_POLY[1023-32* 16 -29])^(crc_i[30]&AHEAD_POLY[1023-32* 16 -30])^(crc_i[31]&AHEAD_POLY[1023-32* 16 -31]);
assign ahead[17] =    (crc_i[0]&AHEAD_POLY[1023-32* 17 ])^(crc_i[1]&AHEAD_POLY[1023-32* 17 -1])^(crc_i[2]&AHEAD_POLY[1023-32*17 -2 ])^(crc_i[3]&AHEAD_POLY[1023-32* 17 -3])^(crc_i[4]&AHEAD_POLY[1023-32* 17 -4])^(crc_i[5]&AHEAD_POLY[1023-32* 17 -5])^(crc_i[6]&AHEAD_POLY[1023-32* 17 -6])^(crc_i[7]&AHEAD_POLY[1023-32* 17 -7])^(crc_i[8]&AHEAD_POLY[1023-32* 17 -8])^(crc_i[9]&AHEAD_POLY[1023-32* 17 -9])^(crc_i[10]&AHEAD_POLY[1023-32* 17 -10])^(crc_i[11]&AHEAD_POLY[1023-32* 17 -11])^(crc_i[12]&AHEAD_POLY[1023-32* 17 -12])^(crc_i[13]&AHEAD_POLY[1023-32* 17 -13])^(crc_i[14]&AHEAD_POLY[1023-32* 17 -14])^(crc_i[15]&AHEAD_POLY[1023-32* 17 -15])^(crc_i[16]&AHEAD_POLY[1023-32* 17 -16])^(crc_i[17]&AHEAD_POLY[1023-32* 17 -17])^(crc_i[18]&AHEAD_POLY[1023-32* 17 -18])^(crc_i[19]&AHEAD_POLY[1023-32* 17 -19])^(crc_i[20]&AHEAD_POLY[1023-32* 17 -20])^(crc_i[21]&AHEAD_POLY[1023-32* 17 -21])^(crc_i[22]&AHEAD_POLY[1023-32* 17 -22])^(crc_i[23]&AHEAD_POLY[1023-32* 17 -23])^(crc_i[24]&AHEAD_POLY[1023-32* 17 -24])^(crc_i[25]&AHEAD_POLY[1023-32* 17 -25])^(crc_i[26]&AHEAD_POLY[1023-32* 17 -26])^(crc_i[27]&AHEAD_POLY[1023-32* 17 -27])^(crc_i[28]&AHEAD_POLY[1023-32* 17 -28])^(crc_i[29]&AHEAD_POLY[1023-32* 17 -29])^(crc_i[30]&AHEAD_POLY[1023-32* 17 -30])^(crc_i[31]&AHEAD_POLY[1023-32* 17 -31]);
assign ahead[18] =    (crc_i[0]&AHEAD_POLY[1023-32* 18 ])^(crc_i[1]&AHEAD_POLY[1023-32* 18 -1])^(crc_i[2]&AHEAD_POLY[1023-32*18 -2 ])^(crc_i[3]&AHEAD_POLY[1023-32* 18 -3])^(crc_i[4]&AHEAD_POLY[1023-32* 18 -4])^(crc_i[5]&AHEAD_POLY[1023-32* 18 -5])^(crc_i[6]&AHEAD_POLY[1023-32* 18 -6])^(crc_i[7]&AHEAD_POLY[1023-32* 18 -7])^(crc_i[8]&AHEAD_POLY[1023-32* 18 -8])^(crc_i[9]&AHEAD_POLY[1023-32* 18 -9])^(crc_i[10]&AHEAD_POLY[1023-32* 18 -10])^(crc_i[11]&AHEAD_POLY[1023-32* 18 -11])^(crc_i[12]&AHEAD_POLY[1023-32* 18 -12])^(crc_i[13]&AHEAD_POLY[1023-32* 18 -13])^(crc_i[14]&AHEAD_POLY[1023-32* 18 -14])^(crc_i[15]&AHEAD_POLY[1023-32* 18 -15])^(crc_i[16]&AHEAD_POLY[1023-32* 18 -16])^(crc_i[17]&AHEAD_POLY[1023-32* 18 -17])^(crc_i[18]&AHEAD_POLY[1023-32* 18 -18])^(crc_i[19]&AHEAD_POLY[1023-32* 18 -19])^(crc_i[20]&AHEAD_POLY[1023-32* 18 -20])^(crc_i[21]&AHEAD_POLY[1023-32* 18 -21])^(crc_i[22]&AHEAD_POLY[1023-32* 18 -22])^(crc_i[23]&AHEAD_POLY[1023-32* 18 -23])^(crc_i[24]&AHEAD_POLY[1023-32* 18 -24])^(crc_i[25]&AHEAD_POLY[1023-32* 18 -25])^(crc_i[26]&AHEAD_POLY[1023-32* 18 -26])^(crc_i[27]&AHEAD_POLY[1023-32* 18 -27])^(crc_i[28]&AHEAD_POLY[1023-32* 18 -28])^(crc_i[29]&AHEAD_POLY[1023-32* 18 -29])^(crc_i[30]&AHEAD_POLY[1023-32* 18 -30])^(crc_i[31]&AHEAD_POLY[1023-32* 18 -31]);
assign ahead[19] =    (crc_i[0]&AHEAD_POLY[1023-32* 19 ])^(crc_i[1]&AHEAD_POLY[1023-32* 19 -1])^(crc_i[2]&AHEAD_POLY[1023-32*19 -2 ])^(crc_i[3]&AHEAD_POLY[1023-32* 19 -3])^(crc_i[4]&AHEAD_POLY[1023-32* 19 -4])^(crc_i[5]&AHEAD_POLY[1023-32* 19 -5])^(crc_i[6]&AHEAD_POLY[1023-32* 19 -6])^(crc_i[7]&AHEAD_POLY[1023-32* 19 -7])^(crc_i[8]&AHEAD_POLY[1023-32* 19 -8])^(crc_i[9]&AHEAD_POLY[1023-32* 19 -9])^(crc_i[10]&AHEAD_POLY[1023-32* 19 -10])^(crc_i[11]&AHEAD_POLY[1023-32* 19 -11])^(crc_i[12]&AHEAD_POLY[1023-32* 19 -12])^(crc_i[13]&AHEAD_POLY[1023-32* 19 -13])^(crc_i[14]&AHEAD_POLY[1023-32* 19 -14])^(crc_i[15]&AHEAD_POLY[1023-32* 19 -15])^(crc_i[16]&AHEAD_POLY[1023-32* 19 -16])^(crc_i[17]&AHEAD_POLY[1023-32* 19 -17])^(crc_i[18]&AHEAD_POLY[1023-32* 19 -18])^(crc_i[19]&AHEAD_POLY[1023-32* 19 -19])^(crc_i[20]&AHEAD_POLY[1023-32* 19 -20])^(crc_i[21]&AHEAD_POLY[1023-32* 19 -21])^(crc_i[22]&AHEAD_POLY[1023-32* 19 -22])^(crc_i[23]&AHEAD_POLY[1023-32* 19 -23])^(crc_i[24]&AHEAD_POLY[1023-32* 19 -24])^(crc_i[25]&AHEAD_POLY[1023-32* 19 -25])^(crc_i[26]&AHEAD_POLY[1023-32* 19 -26])^(crc_i[27]&AHEAD_POLY[1023-32* 19 -27])^(crc_i[28]&AHEAD_POLY[1023-32* 19 -28])^(crc_i[29]&AHEAD_POLY[1023-32* 19 -29])^(crc_i[30]&AHEAD_POLY[1023-32* 19 -30])^(crc_i[31]&AHEAD_POLY[1023-32* 19 -31]);
assign ahead[20] =    (crc_i[0]&AHEAD_POLY[1023-32* 20 ])^(crc_i[1]&AHEAD_POLY[1023-32* 20 -1])^(crc_i[2]&AHEAD_POLY[1023-32*20 -2 ])^(crc_i[3]&AHEAD_POLY[1023-32* 20 -3])^(crc_i[4]&AHEAD_POLY[1023-32* 20 -4])^(crc_i[5]&AHEAD_POLY[1023-32* 20 -5])^(crc_i[6]&AHEAD_POLY[1023-32* 20 -6])^(crc_i[7]&AHEAD_POLY[1023-32* 20 -7])^(crc_i[8]&AHEAD_POLY[1023-32* 20 -8])^(crc_i[9]&AHEAD_POLY[1023-32* 20 -9])^(crc_i[10]&AHEAD_POLY[1023-32* 20 -10])^(crc_i[11]&AHEAD_POLY[1023-32* 20 -11])^(crc_i[12]&AHEAD_POLY[1023-32* 20 -12])^(crc_i[13]&AHEAD_POLY[1023-32* 20 -13])^(crc_i[14]&AHEAD_POLY[1023-32* 20 -14])^(crc_i[15]&AHEAD_POLY[1023-32* 20 -15])^(crc_i[16]&AHEAD_POLY[1023-32* 20 -16])^(crc_i[17]&AHEAD_POLY[1023-32* 20 -17])^(crc_i[18]&AHEAD_POLY[1023-32* 20 -18])^(crc_i[19]&AHEAD_POLY[1023-32* 20 -19])^(crc_i[20]&AHEAD_POLY[1023-32* 20 -20])^(crc_i[21]&AHEAD_POLY[1023-32* 20 -21])^(crc_i[22]&AHEAD_POLY[1023-32* 20 -22])^(crc_i[23]&AHEAD_POLY[1023-32* 20 -23])^(crc_i[24]&AHEAD_POLY[1023-32* 20 -24])^(crc_i[25]&AHEAD_POLY[1023-32* 20 -25])^(crc_i[26]&AHEAD_POLY[1023-32* 20 -26])^(crc_i[27]&AHEAD_POLY[1023-32* 20 -27])^(crc_i[28]&AHEAD_POLY[1023-32* 20 -28])^(crc_i[29]&AHEAD_POLY[1023-32* 20 -29])^(crc_i[30]&AHEAD_POLY[1023-32* 20 -30])^(crc_i[31]&AHEAD_POLY[1023-32* 20 -31]);
assign ahead[21] =    (crc_i[0]&AHEAD_POLY[1023-32* 21 ])^(crc_i[1]&AHEAD_POLY[1023-32* 21 -1])^(crc_i[2]&AHEAD_POLY[1023-32*21 -2 ])^(crc_i[3]&AHEAD_POLY[1023-32* 21 -3])^(crc_i[4]&AHEAD_POLY[1023-32* 21 -4])^(crc_i[5]&AHEAD_POLY[1023-32* 21 -5])^(crc_i[6]&AHEAD_POLY[1023-32* 21 -6])^(crc_i[7]&AHEAD_POLY[1023-32* 21 -7])^(crc_i[8]&AHEAD_POLY[1023-32* 21 -8])^(crc_i[9]&AHEAD_POLY[1023-32* 21 -9])^(crc_i[10]&AHEAD_POLY[1023-32* 21 -10])^(crc_i[11]&AHEAD_POLY[1023-32* 21 -11])^(crc_i[12]&AHEAD_POLY[1023-32* 21 -12])^(crc_i[13]&AHEAD_POLY[1023-32* 21 -13])^(crc_i[14]&AHEAD_POLY[1023-32* 21 -14])^(crc_i[15]&AHEAD_POLY[1023-32* 21 -15])^(crc_i[16]&AHEAD_POLY[1023-32* 21 -16])^(crc_i[17]&AHEAD_POLY[1023-32* 21 -17])^(crc_i[18]&AHEAD_POLY[1023-32* 21 -18])^(crc_i[19]&AHEAD_POLY[1023-32* 21 -19])^(crc_i[20]&AHEAD_POLY[1023-32* 21 -20])^(crc_i[21]&AHEAD_POLY[1023-32* 21 -21])^(crc_i[22]&AHEAD_POLY[1023-32* 21 -22])^(crc_i[23]&AHEAD_POLY[1023-32* 21 -23])^(crc_i[24]&AHEAD_POLY[1023-32* 21 -24])^(crc_i[25]&AHEAD_POLY[1023-32* 21 -25])^(crc_i[26]&AHEAD_POLY[1023-32* 21 -26])^(crc_i[27]&AHEAD_POLY[1023-32* 21 -27])^(crc_i[28]&AHEAD_POLY[1023-32* 21 -28])^(crc_i[29]&AHEAD_POLY[1023-32* 21 -29])^(crc_i[30]&AHEAD_POLY[1023-32* 21 -30])^(crc_i[31]&AHEAD_POLY[1023-32* 21 -31]);
assign ahead[22] =    (crc_i[0]&AHEAD_POLY[1023-32* 22 ])^(crc_i[1]&AHEAD_POLY[1023-32* 22 -1])^(crc_i[2]&AHEAD_POLY[1023-32*22 -2 ])^(crc_i[3]&AHEAD_POLY[1023-32* 22 -3])^(crc_i[4]&AHEAD_POLY[1023-32* 22 -4])^(crc_i[5]&AHEAD_POLY[1023-32* 22 -5])^(crc_i[6]&AHEAD_POLY[1023-32* 22 -6])^(crc_i[7]&AHEAD_POLY[1023-32* 22 -7])^(crc_i[8]&AHEAD_POLY[1023-32* 22 -8])^(crc_i[9]&AHEAD_POLY[1023-32* 22 -9])^(crc_i[10]&AHEAD_POLY[1023-32* 22 -10])^(crc_i[11]&AHEAD_POLY[1023-32* 22 -11])^(crc_i[12]&AHEAD_POLY[1023-32* 22 -12])^(crc_i[13]&AHEAD_POLY[1023-32* 22 -13])^(crc_i[14]&AHEAD_POLY[1023-32* 22 -14])^(crc_i[15]&AHEAD_POLY[1023-32* 22 -15])^(crc_i[16]&AHEAD_POLY[1023-32* 22 -16])^(crc_i[17]&AHEAD_POLY[1023-32* 22 -17])^(crc_i[18]&AHEAD_POLY[1023-32* 22 -18])^(crc_i[19]&AHEAD_POLY[1023-32* 22 -19])^(crc_i[20]&AHEAD_POLY[1023-32* 22 -20])^(crc_i[21]&AHEAD_POLY[1023-32* 22 -21])^(crc_i[22]&AHEAD_POLY[1023-32* 22 -22])^(crc_i[23]&AHEAD_POLY[1023-32* 22 -23])^(crc_i[24]&AHEAD_POLY[1023-32* 22 -24])^(crc_i[25]&AHEAD_POLY[1023-32* 22 -25])^(crc_i[26]&AHEAD_POLY[1023-32* 22 -26])^(crc_i[27]&AHEAD_POLY[1023-32* 22 -27])^(crc_i[28]&AHEAD_POLY[1023-32* 22 -28])^(crc_i[29]&AHEAD_POLY[1023-32* 22 -29])^(crc_i[30]&AHEAD_POLY[1023-32* 22 -30])^(crc_i[31]&AHEAD_POLY[1023-32* 22 -31]);
assign ahead[23] =    (crc_i[0]&AHEAD_POLY[1023-32* 23 ])^(crc_i[1]&AHEAD_POLY[1023-32* 23 -1])^(crc_i[2]&AHEAD_POLY[1023-32*23 -2 ])^(crc_i[3]&AHEAD_POLY[1023-32* 23 -3])^(crc_i[4]&AHEAD_POLY[1023-32* 23 -4])^(crc_i[5]&AHEAD_POLY[1023-32* 23 -5])^(crc_i[6]&AHEAD_POLY[1023-32* 23 -6])^(crc_i[7]&AHEAD_POLY[1023-32* 23 -7])^(crc_i[8]&AHEAD_POLY[1023-32* 23 -8])^(crc_i[9]&AHEAD_POLY[1023-32* 23 -9])^(crc_i[10]&AHEAD_POLY[1023-32* 23 -10])^(crc_i[11]&AHEAD_POLY[1023-32* 23 -11])^(crc_i[12]&AHEAD_POLY[1023-32* 23 -12])^(crc_i[13]&AHEAD_POLY[1023-32* 23 -13])^(crc_i[14]&AHEAD_POLY[1023-32* 23 -14])^(crc_i[15]&AHEAD_POLY[1023-32* 23 -15])^(crc_i[16]&AHEAD_POLY[1023-32* 23 -16])^(crc_i[17]&AHEAD_POLY[1023-32* 23 -17])^(crc_i[18]&AHEAD_POLY[1023-32* 23 -18])^(crc_i[19]&AHEAD_POLY[1023-32* 23 -19])^(crc_i[20]&AHEAD_POLY[1023-32* 23 -20])^(crc_i[21]&AHEAD_POLY[1023-32* 23 -21])^(crc_i[22]&AHEAD_POLY[1023-32* 23 -22])^(crc_i[23]&AHEAD_POLY[1023-32* 23 -23])^(crc_i[24]&AHEAD_POLY[1023-32* 23 -24])^(crc_i[25]&AHEAD_POLY[1023-32* 23 -25])^(crc_i[26]&AHEAD_POLY[1023-32* 23 -26])^(crc_i[27]&AHEAD_POLY[1023-32* 23 -27])^(crc_i[28]&AHEAD_POLY[1023-32* 23 -28])^(crc_i[29]&AHEAD_POLY[1023-32* 23 -29])^(crc_i[30]&AHEAD_POLY[1023-32* 23 -30])^(crc_i[31]&AHEAD_POLY[1023-32* 23 -31]);
assign ahead[24] =    (crc_i[0]&AHEAD_POLY[1023-32* 24 ])^(crc_i[1]&AHEAD_POLY[1023-32* 24 -1])^(crc_i[2]&AHEAD_POLY[1023-32*24 -2 ])^(crc_i[3]&AHEAD_POLY[1023-32* 24 -3])^(crc_i[4]&AHEAD_POLY[1023-32* 24 -4])^(crc_i[5]&AHEAD_POLY[1023-32* 24 -5])^(crc_i[6]&AHEAD_POLY[1023-32* 24 -6])^(crc_i[7]&AHEAD_POLY[1023-32* 24 -7])^(crc_i[8]&AHEAD_POLY[1023-32* 24 -8])^(crc_i[9]&AHEAD_POLY[1023-32* 24 -9])^(crc_i[10]&AHEAD_POLY[1023-32* 24 -10])^(crc_i[11]&AHEAD_POLY[1023-32* 24 -11])^(crc_i[12]&AHEAD_POLY[1023-32* 24 -12])^(crc_i[13]&AHEAD_POLY[1023-32* 24 -13])^(crc_i[14]&AHEAD_POLY[1023-32* 24 -14])^(crc_i[15]&AHEAD_POLY[1023-32* 24 -15])^(crc_i[16]&AHEAD_POLY[1023-32* 24 -16])^(crc_i[17]&AHEAD_POLY[1023-32* 24 -17])^(crc_i[18]&AHEAD_POLY[1023-32* 24 -18])^(crc_i[19]&AHEAD_POLY[1023-32* 24 -19])^(crc_i[20]&AHEAD_POLY[1023-32* 24 -20])^(crc_i[21]&AHEAD_POLY[1023-32* 24 -21])^(crc_i[22]&AHEAD_POLY[1023-32* 24 -22])^(crc_i[23]&AHEAD_POLY[1023-32* 24 -23])^(crc_i[24]&AHEAD_POLY[1023-32* 24 -24])^(crc_i[25]&AHEAD_POLY[1023-32* 24 -25])^(crc_i[26]&AHEAD_POLY[1023-32* 24 -26])^(crc_i[27]&AHEAD_POLY[1023-32* 24 -27])^(crc_i[28]&AHEAD_POLY[1023-32* 24 -28])^(crc_i[29]&AHEAD_POLY[1023-32* 24 -29])^(crc_i[30]&AHEAD_POLY[1023-32* 24 -30])^(crc_i[31]&AHEAD_POLY[1023-32* 24 -31]);
assign ahead[25] =    (crc_i[0]&AHEAD_POLY[1023-32* 25 ])^(crc_i[1]&AHEAD_POLY[1023-32* 25 -1])^(crc_i[2]&AHEAD_POLY[1023-32*25 -2 ])^(crc_i[3]&AHEAD_POLY[1023-32* 25 -3])^(crc_i[4]&AHEAD_POLY[1023-32* 25 -4])^(crc_i[5]&AHEAD_POLY[1023-32* 25 -5])^(crc_i[6]&AHEAD_POLY[1023-32* 25 -6])^(crc_i[7]&AHEAD_POLY[1023-32* 25 -7])^(crc_i[8]&AHEAD_POLY[1023-32* 25 -8])^(crc_i[9]&AHEAD_POLY[1023-32* 25 -9])^(crc_i[10]&AHEAD_POLY[1023-32* 25 -10])^(crc_i[11]&AHEAD_POLY[1023-32* 25 -11])^(crc_i[12]&AHEAD_POLY[1023-32* 25 -12])^(crc_i[13]&AHEAD_POLY[1023-32* 25 -13])^(crc_i[14]&AHEAD_POLY[1023-32* 25 -14])^(crc_i[15]&AHEAD_POLY[1023-32* 25 -15])^(crc_i[16]&AHEAD_POLY[1023-32* 25 -16])^(crc_i[17]&AHEAD_POLY[1023-32* 25 -17])^(crc_i[18]&AHEAD_POLY[1023-32* 25 -18])^(crc_i[19]&AHEAD_POLY[1023-32* 25 -19])^(crc_i[20]&AHEAD_POLY[1023-32* 25 -20])^(crc_i[21]&AHEAD_POLY[1023-32* 25 -21])^(crc_i[22]&AHEAD_POLY[1023-32* 25 -22])^(crc_i[23]&AHEAD_POLY[1023-32* 25 -23])^(crc_i[24]&AHEAD_POLY[1023-32* 25 -24])^(crc_i[25]&AHEAD_POLY[1023-32* 25 -25])^(crc_i[26]&AHEAD_POLY[1023-32* 25 -26])^(crc_i[27]&AHEAD_POLY[1023-32* 25 -27])^(crc_i[28]&AHEAD_POLY[1023-32* 25 -28])^(crc_i[29]&AHEAD_POLY[1023-32* 25 -29])^(crc_i[30]&AHEAD_POLY[1023-32* 25 -30])^(crc_i[31]&AHEAD_POLY[1023-32* 25 -31]);
assign ahead[26] =    (crc_i[0]&AHEAD_POLY[1023-32* 26 ])^(crc_i[1]&AHEAD_POLY[1023-32* 26 -1])^(crc_i[2]&AHEAD_POLY[1023-32*26 -2 ])^(crc_i[3]&AHEAD_POLY[1023-32* 26 -3])^(crc_i[4]&AHEAD_POLY[1023-32* 26 -4])^(crc_i[5]&AHEAD_POLY[1023-32* 26 -5])^(crc_i[6]&AHEAD_POLY[1023-32* 26 -6])^(crc_i[7]&AHEAD_POLY[1023-32* 26 -7])^(crc_i[8]&AHEAD_POLY[1023-32* 26 -8])^(crc_i[9]&AHEAD_POLY[1023-32* 26 -9])^(crc_i[10]&AHEAD_POLY[1023-32* 26 -10])^(crc_i[11]&AHEAD_POLY[1023-32* 26 -11])^(crc_i[12]&AHEAD_POLY[1023-32* 26 -12])^(crc_i[13]&AHEAD_POLY[1023-32* 26 -13])^(crc_i[14]&AHEAD_POLY[1023-32* 26 -14])^(crc_i[15]&AHEAD_POLY[1023-32* 26 -15])^(crc_i[16]&AHEAD_POLY[1023-32* 26 -16])^(crc_i[17]&AHEAD_POLY[1023-32* 26 -17])^(crc_i[18]&AHEAD_POLY[1023-32* 26 -18])^(crc_i[19]&AHEAD_POLY[1023-32* 26 -19])^(crc_i[20]&AHEAD_POLY[1023-32* 26 -20])^(crc_i[21]&AHEAD_POLY[1023-32* 26 -21])^(crc_i[22]&AHEAD_POLY[1023-32* 26 -22])^(crc_i[23]&AHEAD_POLY[1023-32* 26 -23])^(crc_i[24]&AHEAD_POLY[1023-32* 26 -24])^(crc_i[25]&AHEAD_POLY[1023-32* 26 -25])^(crc_i[26]&AHEAD_POLY[1023-32* 26 -26])^(crc_i[27]&AHEAD_POLY[1023-32* 26 -27])^(crc_i[28]&AHEAD_POLY[1023-32* 26 -28])^(crc_i[29]&AHEAD_POLY[1023-32* 26 -29])^(crc_i[30]&AHEAD_POLY[1023-32* 26 -30])^(crc_i[31]&AHEAD_POLY[1023-32* 26 -31]);
assign ahead[27] =    (crc_i[0]&AHEAD_POLY[1023-32* 27 ])^(crc_i[1]&AHEAD_POLY[1023-32* 27 -1])^(crc_i[2]&AHEAD_POLY[1023-32*27 -2 ])^(crc_i[3]&AHEAD_POLY[1023-32* 27 -3])^(crc_i[4]&AHEAD_POLY[1023-32* 27 -4])^(crc_i[5]&AHEAD_POLY[1023-32* 27 -5])^(crc_i[6]&AHEAD_POLY[1023-32* 27 -6])^(crc_i[7]&AHEAD_POLY[1023-32* 27 -7])^(crc_i[8]&AHEAD_POLY[1023-32* 27 -8])^(crc_i[9]&AHEAD_POLY[1023-32* 27 -9])^(crc_i[10]&AHEAD_POLY[1023-32* 27 -10])^(crc_i[11]&AHEAD_POLY[1023-32* 27 -11])^(crc_i[12]&AHEAD_POLY[1023-32* 27 -12])^(crc_i[13]&AHEAD_POLY[1023-32* 27 -13])^(crc_i[14]&AHEAD_POLY[1023-32* 27 -14])^(crc_i[15]&AHEAD_POLY[1023-32* 27 -15])^(crc_i[16]&AHEAD_POLY[1023-32* 27 -16])^(crc_i[17]&AHEAD_POLY[1023-32* 27 -17])^(crc_i[18]&AHEAD_POLY[1023-32* 27 -18])^(crc_i[19]&AHEAD_POLY[1023-32* 27 -19])^(crc_i[20]&AHEAD_POLY[1023-32* 27 -20])^(crc_i[21]&AHEAD_POLY[1023-32* 27 -21])^(crc_i[22]&AHEAD_POLY[1023-32* 27 -22])^(crc_i[23]&AHEAD_POLY[1023-32* 27 -23])^(crc_i[24]&AHEAD_POLY[1023-32* 27 -24])^(crc_i[25]&AHEAD_POLY[1023-32* 27 -25])^(crc_i[26]&AHEAD_POLY[1023-32* 27 -26])^(crc_i[27]&AHEAD_POLY[1023-32* 27 -27])^(crc_i[28]&AHEAD_POLY[1023-32* 27 -28])^(crc_i[29]&AHEAD_POLY[1023-32* 27 -29])^(crc_i[30]&AHEAD_POLY[1023-32* 27 -30])^(crc_i[31]&AHEAD_POLY[1023-32* 27 -31]);
assign ahead[28] =    (crc_i[0]&AHEAD_POLY[1023-32* 28 ])^(crc_i[1]&AHEAD_POLY[1023-32* 28 -1])^(crc_i[2]&AHEAD_POLY[1023-32*28 -2 ])^(crc_i[3]&AHEAD_POLY[1023-32* 28 -3])^(crc_i[4]&AHEAD_POLY[1023-32* 28 -4])^(crc_i[5]&AHEAD_POLY[1023-32* 28 -5])^(crc_i[6]&AHEAD_POLY[1023-32* 28 -6])^(crc_i[7]&AHEAD_POLY[1023-32* 28 -7])^(crc_i[8]&AHEAD_POLY[1023-32* 28 -8])^(crc_i[9]&AHEAD_POLY[1023-32* 28 -9])^(crc_i[10]&AHEAD_POLY[1023-32* 28 -10])^(crc_i[11]&AHEAD_POLY[1023-32* 28 -11])^(crc_i[12]&AHEAD_POLY[1023-32* 28 -12])^(crc_i[13]&AHEAD_POLY[1023-32* 28 -13])^(crc_i[14]&AHEAD_POLY[1023-32* 28 -14])^(crc_i[15]&AHEAD_POLY[1023-32* 28 -15])^(crc_i[16]&AHEAD_POLY[1023-32* 28 -16])^(crc_i[17]&AHEAD_POLY[1023-32* 28 -17])^(crc_i[18]&AHEAD_POLY[1023-32* 28 -18])^(crc_i[19]&AHEAD_POLY[1023-32* 28 -19])^(crc_i[20]&AHEAD_POLY[1023-32* 28 -20])^(crc_i[21]&AHEAD_POLY[1023-32* 28 -21])^(crc_i[22]&AHEAD_POLY[1023-32* 28 -22])^(crc_i[23]&AHEAD_POLY[1023-32* 28 -23])^(crc_i[24]&AHEAD_POLY[1023-32* 28 -24])^(crc_i[25]&AHEAD_POLY[1023-32* 28 -25])^(crc_i[26]&AHEAD_POLY[1023-32* 28 -26])^(crc_i[27]&AHEAD_POLY[1023-32* 28 -27])^(crc_i[28]&AHEAD_POLY[1023-32* 28 -28])^(crc_i[29]&AHEAD_POLY[1023-32* 28 -29])^(crc_i[30]&AHEAD_POLY[1023-32* 28 -30])^(crc_i[31]&AHEAD_POLY[1023-32* 28 -31]);
assign ahead[29] =    (crc_i[0]&AHEAD_POLY[1023-32* 29 ])^(crc_i[1]&AHEAD_POLY[1023-32* 29 -1])^(crc_i[2]&AHEAD_POLY[1023-32*29 -2 ])^(crc_i[3]&AHEAD_POLY[1023-32* 29 -3])^(crc_i[4]&AHEAD_POLY[1023-32* 29 -4])^(crc_i[5]&AHEAD_POLY[1023-32* 29 -5])^(crc_i[6]&AHEAD_POLY[1023-32* 29 -6])^(crc_i[7]&AHEAD_POLY[1023-32* 29 -7])^(crc_i[8]&AHEAD_POLY[1023-32* 29 -8])^(crc_i[9]&AHEAD_POLY[1023-32* 29 -9])^(crc_i[10]&AHEAD_POLY[1023-32* 29 -10])^(crc_i[11]&AHEAD_POLY[1023-32* 29 -11])^(crc_i[12]&AHEAD_POLY[1023-32* 29 -12])^(crc_i[13]&AHEAD_POLY[1023-32* 29 -13])^(crc_i[14]&AHEAD_POLY[1023-32* 29 -14])^(crc_i[15]&AHEAD_POLY[1023-32* 29 -15])^(crc_i[16]&AHEAD_POLY[1023-32* 29 -16])^(crc_i[17]&AHEAD_POLY[1023-32* 29 -17])^(crc_i[18]&AHEAD_POLY[1023-32* 29 -18])^(crc_i[19]&AHEAD_POLY[1023-32* 29 -19])^(crc_i[20]&AHEAD_POLY[1023-32* 29 -20])^(crc_i[21]&AHEAD_POLY[1023-32* 29 -21])^(crc_i[22]&AHEAD_POLY[1023-32* 29 -22])^(crc_i[23]&AHEAD_POLY[1023-32* 29 -23])^(crc_i[24]&AHEAD_POLY[1023-32* 29 -24])^(crc_i[25]&AHEAD_POLY[1023-32* 29 -25])^(crc_i[26]&AHEAD_POLY[1023-32* 29 -26])^(crc_i[27]&AHEAD_POLY[1023-32* 29 -27])^(crc_i[28]&AHEAD_POLY[1023-32* 29 -28])^(crc_i[29]&AHEAD_POLY[1023-32* 29 -29])^(crc_i[30]&AHEAD_POLY[1023-32* 29 -30])^(crc_i[31]&AHEAD_POLY[1023-32* 29 -31]);
assign ahead[30] =    (crc_i[0]&AHEAD_POLY[1023-32* 30 ])^(crc_i[1]&AHEAD_POLY[1023-32* 30 -1])^(crc_i[2]&AHEAD_POLY[1023-32*30 -2 ])^(crc_i[3]&AHEAD_POLY[1023-32* 30 -3])^(crc_i[4]&AHEAD_POLY[1023-32* 30 -4])^(crc_i[5]&AHEAD_POLY[1023-32* 30 -5])^(crc_i[6]&AHEAD_POLY[1023-32* 30 -6])^(crc_i[7]&AHEAD_POLY[1023-32* 30 -7])^(crc_i[8]&AHEAD_POLY[1023-32* 30 -8])^(crc_i[9]&AHEAD_POLY[1023-32* 30 -9])^(crc_i[10]&AHEAD_POLY[1023-32* 30 -10])^(crc_i[11]&AHEAD_POLY[1023-32* 30 -11])^(crc_i[12]&AHEAD_POLY[1023-32* 30 -12])^(crc_i[13]&AHEAD_POLY[1023-32* 30 -13])^(crc_i[14]&AHEAD_POLY[1023-32* 30 -14])^(crc_i[15]&AHEAD_POLY[1023-32* 30 -15])^(crc_i[16]&AHEAD_POLY[1023-32* 30 -16])^(crc_i[17]&AHEAD_POLY[1023-32* 30 -17])^(crc_i[18]&AHEAD_POLY[1023-32* 30 -18])^(crc_i[19]&AHEAD_POLY[1023-32* 30 -19])^(crc_i[20]&AHEAD_POLY[1023-32* 30 -20])^(crc_i[21]&AHEAD_POLY[1023-32* 30 -21])^(crc_i[22]&AHEAD_POLY[1023-32* 30 -22])^(crc_i[23]&AHEAD_POLY[1023-32* 30 -23])^(crc_i[24]&AHEAD_POLY[1023-32* 30 -24])^(crc_i[25]&AHEAD_POLY[1023-32* 30 -25])^(crc_i[26]&AHEAD_POLY[1023-32* 30 -26])^(crc_i[27]&AHEAD_POLY[1023-32* 30 -27])^(crc_i[28]&AHEAD_POLY[1023-32* 30 -28])^(crc_i[29]&AHEAD_POLY[1023-32* 30 -29])^(crc_i[30]&AHEAD_POLY[1023-32* 30 -30])^(crc_i[31]&AHEAD_POLY[1023-32* 30 -31]);
assign ahead[31] =    (crc_i[0]&AHEAD_POLY[1023-32* 31 ])^(crc_i[1]&AHEAD_POLY[1023-32* 31 -1])^(crc_i[2]&AHEAD_POLY[1023-32*31 -2 ])^(crc_i[3]&AHEAD_POLY[1023-32* 31 -3])^(crc_i[4]&AHEAD_POLY[1023-32* 31 -4])^(crc_i[5]&AHEAD_POLY[1023-32* 31 -5])^(crc_i[6]&AHEAD_POLY[1023-32* 31 -6])^(crc_i[7]&AHEAD_POLY[1023-32* 31 -7])^(crc_i[8]&AHEAD_POLY[1023-32* 31 -8])^(crc_i[9]&AHEAD_POLY[1023-32* 31 -9])^(crc_i[10]&AHEAD_POLY[1023-32* 31 -10])^(crc_i[11]&AHEAD_POLY[1023-32* 31 -11])^(crc_i[12]&AHEAD_POLY[1023-32* 31 -12])^(crc_i[13]&AHEAD_POLY[1023-32* 31 -13])^(crc_i[14]&AHEAD_POLY[1023-32* 31 -14])^(crc_i[15]&AHEAD_POLY[1023-32* 31 -15])^(crc_i[16]&AHEAD_POLY[1023-32* 31 -16])^(crc_i[17]&AHEAD_POLY[1023-32* 31 -17])^(crc_i[18]&AHEAD_POLY[1023-32* 31 -18])^(crc_i[19]&AHEAD_POLY[1023-32* 31 -19])^(crc_i[20]&AHEAD_POLY[1023-32* 31 -20])^(crc_i[21]&AHEAD_POLY[1023-32* 31 -21])^(crc_i[22]&AHEAD_POLY[1023-32* 31 -22])^(crc_i[23]&AHEAD_POLY[1023-32* 31 -23])^(crc_i[24]&AHEAD_POLY[1023-32* 31 -24])^(crc_i[25]&AHEAD_POLY[1023-32* 31 -25])^(crc_i[26]&AHEAD_POLY[1023-32* 31 -26])^(crc_i[27]&AHEAD_POLY[1023-32* 31 -27])^(crc_i[28]&AHEAD_POLY[1023-32* 31 -28])^(crc_i[29]&AHEAD_POLY[1023-32* 31 -29])^(crc_i[30]&AHEAD_POLY[1023-32* 31 -30])^(crc_i[31]&AHEAD_POLY[1023-32* 31 -31]);

























// assign crc_en_o = crc_en_i ;
// assign crc_o = CRC32_ahead(crc_i) ;

always @(posedge clk  ) begin
    // if (rst) begin
    //     // reset
    //     crc_en_o    <= 'b0 ;
    //     crc_o       <= 'b0 ;
    // end
    // else begin
        crc_en_o <= crc_en_i     ;
        crc_o    <= ahead        ;
    // end
end



//*********************
endmodule   