


module layer_1_new 
    # ( parameter  LUT_NUM_ONE_EQUATION    		= 171 ,      // and thre are 32 equation
    			   LUT_OUT_NUM_ONE_EQUATION     = 174 ,                   
    	           BUS_WIDTH  		            = LUT_NUM_ONE_EQUATION*5  
        )
( 
            input	            		clk      ,   
            input	            		rst      ,   
            input      [BUS_WIDTH-1:0]    	din      ,
            output reg [LUT_OUT_NUM_ONE_EQUATION*32-1:0]       dout 				      

 ) ;






parameter  [0:LUT_NUM_ONE_EQUATION*64*16-1] POLY  = { 
64'haaaaaaaa5555aaaa,
64'h3333cccc55aa55aa,
64'h5a5a5a5a0ff00ff0,
64'hcccccccc0f0ff0f0,
64'hffff0000c3c33c3c,
64'h669999663333cccc,
64'h696996965a5a5a5a,
64'hf0f0f0f05a5a5a5a,
64'hffff0000ffff0000,
64'ha55aa55ac33cc33c,
64'haa5555aacccccccc,
64'h55aa55aa3c3c3c3c,
64'h9966996600000000,
64'h6996699633cc33cc,
64'h0ff00ff000000000,
64'hffff0000a55aa55a,
64'h3cc3c33cf00f0ff0,
64'h5a5a5a5ac3c33c3c,
64'hffff000099996666,
64'h966969960f0ff0f0,
64'hcc3333cc5aa5a55a,
64'hcccccccc5555aaaa,
64'h6699996696969696,
64'h3cc3c33c66999966,
64'hff00ff0099996666,
64'h699669960ff00ff0,
64'h0f0ff0f03333cccc,
64'h9696969699669966,
64'h00ffff0066999966,
64'hffff0000aaaaaaaa,
64'hcccccccc33cc33cc,
64'h9966996696969696,
64'h3c3c3c3caaaaaaaa,
64'hc3c33c3cf0f0f0f0,
64'h96969696aa5555aa,
64'h00000000ffff0000,
64'h0ff00ff03cc3c33c,
64'h33cc33cc99996666,
64'h9669699655aa55aa,
64'hf00f0ff03333cccc,
64'hc33cc33c5a5a5a5a,
64'hf00f0ff0a5a55a5a,
64'ha5a55a5a3c3c3c3c,
64'hcccccccccc3333cc,
64'hffff000069966996,
64'hc33cc33c0ff00ff0,
64'h5555aaaa69966996,
64'hf0f0f0f0f00f0ff0,
64'hff00ff00ff00ff00,
64'hff00ff0069699696,
64'hf0f0f0f0aaaaaaaa,
64'ha5a55a5a00000000,
64'h3333ccccaa5555aa,
64'haa5555aaff00ff00,
64'h00ffff005555aaaa,
64'hc3c33c3ccccccccc,
64'hff00ff00c3c33c3c,
64'hc33cc33cc33cc33c,
64'ha5a55a5a5a5a5a5a,
64'h966969963cc3c33c,
64'ha55aa55a69966996,
64'h5555aaaa5a5a5a5a,
64'h5a5a5a5a00000000,
64'h5aa5a55a3333cccc,
64'h9696969699996666,
64'h0ff00ff00f0ff0f0,
64'h00ffff00aaaaaaaa,
64'h5aa5a55a69966996,
64'hc3c33c3c69966996,
64'h5aa5a55af00f0ff0,
64'hff00ff00ff00ff00,
64'hf00f0ff05a5a5a5a,
64'h0ff00ff0cc3333cc,
64'hcc3333cc0f0ff0f0,
64'h0f0ff0f0cccccccc,
64'h33cc33cc00ffff00,
64'hcccccccc3cc3c33c,
64'hc33cc33cc3c33c3c,
64'h699669960ff00ff0,
64'hcc3333cc66666666,
64'h5555aaaaffff0000,
64'h5aa5a55a69966996,
64'h0f0ff0f096696996,
64'hcc3333cc66666666,
64'h0f0ff0f066999966,
64'h000000000f0ff0f0,
64'h00ffff00c33cc33c,
64'h3c3c3c3cc3c33c3c,
64'hffff000099996666,
64'h00ffff00ffff0000,
64'h5a5a5a5a0f0ff0f0,
64'hff00ff005aa5a55a,
64'hc3c33c3c00000000,
64'h55aa55aacccccccc,
64'h5a5a5a5a0f0ff0f0,
64'hc3c33c3c5555aaaa,
64'h699669960ff00ff0,
64'hcc3333cc3333cccc,
64'h9669699600ffff00,
64'haaaaaaaa69699696,
64'h96969696c3c33c3c,
64'hc33cc33c69699696,
64'h6969969600000000,
64'hcc3333cc33cc33cc,
64'h3c3c3c3c0ff00ff0,
64'h66999966a5a55a5a,
64'h69699696aa5555aa,
64'h5555aaaa99996666,
64'h5a5a5a5aaa5555aa,
64'h5555aaaa96696996,
64'h3333cccc5a5a5a5a,
64'h6996699696969696,
64'h996699665aa5a55a,
64'h5a5a5a5ac33cc33c,
64'hcc3333cc0f0ff0f0,
64'h55aa55aa3cc3c33c,
64'h55aa55aa5a5a5a5a,
64'h969696965555aaaa,
64'hc33cc33c99996666,
64'h9999666600ffff00,
64'h5aa5a55a99996666,
64'hc3c33c3c5a5a5a5a,
64'h6996699669699696,
64'ha5a55a5a33cc33cc,
64'haa5555aaaaaaaaaa,
64'h3333cccc66999966,
64'h5a5a5a5aaaaaaaaa,
64'hcccccccc99996666,
64'ha5a55a5acccccccc,
64'hcc3333ccc3c33c3c,
64'h0ff00ff000ffff00,
64'h9966996655aa55aa,
64'h000000005aa5a55a,
64'h96696996ffff0000,
64'h5aa5a55a3333cccc,
64'haaaaaaaa66999966,
64'haaaaaaaaffff0000,
64'hc3c33c3c5555aaaa,
64'hcc3333cc69966996,
64'h55aa55aa3333cccc,
64'h69699696f0f0f0f0,
64'h0ff00ff0c3c33c3c,
64'haaaaaaaa5555aaaa,
64'h5555aaaa3c3c3c3c,
64'h96696996ff00ff00,
64'ha5a55a5a66999966,
64'h3c3c3c3cff00ff00,
64'hccccccccc3c33c3c,
64'h696996965555aaaa,
64'h0ff00ff099996666,
64'h55aa55aaaaaaaaaa,
64'h9966996600000000,
64'h0ff00ff0c33cc33c,
64'ha5a55a5af0f0f0f0,
64'hffff000055aa55aa,
64'hcccccccc55aa55aa,
64'ha5a55a5a55aa55aa,
64'h99669966aaaaaaaa,
64'h33cc33ccf00f0ff0,
64'hff00ff0000ffff00,
64'h5aa5a55a3333cccc,
64'h3cc3c33c66666666,
64'h96696996aa5555aa,
64'h6699996699669966,
64'hffff0000a55aa55a,
64'h5a5a5a5a00000000,
64'h0f0ff0f069966996,
64'ha5a55a5af0f0f0f0,
64'h5a5a5a5acccccccc,
64'hcc3333cccc3333cc,
64'h66999966cccccccc,
64'h0f0ff0f03c3c3c3c,
64'h996699660ff00ff0,
64'hf00f0ff0aa5555aa,
64'hcc3333cc55aa55aa,
64'h96696996f0f0f0f0,
64'h33cc33cc3333cccc,
64'hc3c33c3c3c3c3c3c,
64'h996699660ff00ff0,
64'h3cc3c33cc33cc33c,
64'h96696996a55aa55a,
64'h3c3c3c3ca5a55a5a,
64'haaaaaaaaf00f0ff0,
64'ha55aa55a5aa5a55a,
64'haaaaaaaa3c3c3c3c,
64'h0000000066666666,
64'hcc3333ccf00f0ff0,
64'haa5555aaaa5555aa,
64'h3333cccc66999966,
64'hff00ff0099669966,
64'haa5555aa5555aaaa,
64'haa5555aa5aa5a55a,
64'haaaaaaaa96696996,
64'hf0f0f0f069699696,
64'h3333ccccc33cc33c,
64'h5aa5a55a66999966,
64'h96696996ffff0000,
64'haaaaaaaa5aa5a55a,
64'ha5a55a5a69966996,
64'hcc3333cc0ff00ff0,
64'h5555aaaaffff0000,
64'h66999966ff00ff00,
64'h3c3c3c3ca5a55a5a,
64'h6699996699669966,
64'hcccccccc69966996,
64'h66666666cccccccc,
64'hc3c33c3c99996666,
64'hc33cc33c00ffff00,
64'h3c3c3c3cff00ff00,
64'hffff0000a55aa55a,
64'h0ff00ff05a5a5a5a,
64'h00ffff0099669966,
64'ha55aa55a33cc33cc,
64'hffff000000000000,
64'hc3c33c3c5aa5a55a,
64'h99669966f0f0f0f0,
64'hcc3333cc0ff00ff0,
64'h5aa5a55a00000000,
64'h5555aaaa0f0ff0f0,
64'h0f0ff0f000000000,
64'hffff0000cc3333cc,
64'h6666666600ffff00,
64'hc33cc33ca55aa55a,
64'hffff000096969696,
64'h0000000055aa55aa,
64'h6996699666999966,
64'h9696969666666666,
64'ha55aa55a69966996,
64'h66666666c3c33c3c,
64'haa5555aa96969696,
64'h5555aaaaaa5555aa,
64'hf00f0ff0f0f0f0f0,
64'hff00ff0069699696,
64'hff00ff00c3c33c3c,
64'h5555aaaa66666666,
64'h969696960f0ff0f0,
64'h5aa5a55ac33cc33c,
64'h33cc33cccccccccc,
64'hcc3333ccff00ff00,
64'hff00ff003333cccc,
64'h00000000aaaaaaaa,
64'h0f0ff0f05aa5a55a,
64'h3cc3c33c96969696,
64'haaaaaaaa99996666,
64'h5a5a5a5af0f0f0f0,
64'h9999666699669966,
64'hf0f0f0f033cc33cc,
64'h3cc3c33ca55aa55a,
64'h969696960f0ff0f0,
64'hffff000096696996,
64'h9999666600ffff00,
64'h999966663cc3c33c,
64'ha55aa55a00ffff00,
64'h00ffff005555aaaa,
64'h00ffff00c33cc33c,
64'h0ff00ff066666666,
64'h9669699600000000,
64'h696996963333cccc,
64'h33cc33cc5555aaaa,
64'h55aa55aacccccccc,
64'h669999665a5a5a5a,
64'haa5555aa0ff00ff0,
64'h3333cccc5aa5a55a,
64'h9669699633cc33cc,
64'h00000000f00f0ff0,
64'hc3c33c3c96696996,
64'h9999666633cc33cc,
64'hc33cc33c00000000,
64'h96969696f0f0f0f0,
64'hff00ff0096969696,
64'h0f0ff0f055aa55aa,
64'hff00ff0066666666,
64'h3c3c3c3c3cc3c33c,
64'h669999663cc3c33c,
64'h3c3c3c3c00ffff00,
64'haa5555aa5555aaaa,
64'hf0f0f0f033cc33cc,
64'ha5a55a5a0f0ff0f0,
64'hc33cc33c55aa55aa,
64'h5aa5a55a5a5a5a5a,
64'h96696996ffff0000,
64'h3c3c3c3c5aa5a55a,
64'h3333cccca55aa55a,
64'h5555aaaaaa5555aa,
64'hc33cc33c3c3c3c3c,
64'h3333cccc00000000,
64'h3c3c3c3c96696996,
64'h5aa5a55a3cc3c33c,
64'h6996699696969696,
64'h5aa5a55ac3c33c3c,
64'haaaaaaaa55aa55aa,
64'hff00ff005aa5a55a,
64'h996699660ff00ff0,
64'hffff000096969696,
64'h55aa55aaaaaaaaaa,
64'hc33cc33c55aa55aa,
64'h00ffff0066999966,
64'hcc3333ccaaaaaaaa,
64'hcc3333ccf0f0f0f0,
64'h69966996ff00ff00,
64'hcc3333cc66666666,
64'hffff0000aa5555aa,
64'hc33cc33cf0f0f0f0,
64'h000000005555aaaa,
64'hcccccccc69966996,
64'h55aa55aaa55aa55a,
64'h3333cccc69966996,
64'haa5555aaaaaaaaaa,
64'h699669960f0ff0f0,
64'h9966996600ffff00,
64'ha55aa55a33cc33cc,
64'h00ffff0099996666,
64'h3333cccc96969696,
64'hc33cc33c99996666,
64'h9999666696696996,
64'h6969969699669966,
64'hffff0000c33cc33c,
64'h5aa5a55acc3333cc,
64'h699669965aa5a55a,
64'hc33cc33cff00ff00,
64'hcc3333cc5aa5a55a,
64'h6699996699669966,
64'h55aa55aacccccccc,
64'h3333cccc96969696,
64'ha5a55a5a5555aaaa,
64'h3c3c3c3c96969696,
64'h6699996699669966,
64'hffff0000c33cc33c,
64'h96696996a5a55a5a,
64'h33cc33cccccccccc,
64'h69699696c3c33c3c,
64'hc33cc33c66666666,
64'h3c3c3c3c3c3c3c3c,
64'h966969965a5a5a5a,
64'h699669960ff00ff0,
64'ha5a55a5a5555aaaa,
64'h5aa5a55a99996666,
64'h00000000cc3333cc,
64'haaaaaaaaaaaaaaaa,
64'h3c3c3c3c5a5a5a5a,
64'hcccccccc69699696,
64'h66666666aaaaaaaa,
64'hcc3333cc66666666,
64'h6996699696696996,
64'hcc3333ccf0f0f0f0,
64'haa5555aa55aa55aa,
64'ha5a55a5a0ff00ff0,
64'h6666666666666666,
64'h99996666a55aa55a,
64'h00000000ffff0000,
64'h3cc3c33cc3c33c3c,
64'h996699665555aaaa,
64'h3c3c3c3c0ff00ff0,
64'haa5555aa66666666,
64'ha5a55a5a96969696,
64'h6699996666666666,
64'h5aa5a55a00000000,
64'h0f0ff0f0f00f0ff0,
64'h96696996ff00ff00,
64'h5555aaaa3333cccc,
64'h969696963333cccc,
64'h966969963333cccc,
64'hf00f0ff0cccccccc,
64'h3cc3c33c00ffff00,
64'h00ffff005555aaaa,
64'h969696965a5a5a5a,
64'h6666666696969696,
64'h000000003333cccc,
64'h0ff00ff069699696,
64'h5555aaaacc3333cc,
64'hc33cc33c00000000,
64'hf00f0ff03cc3c33c,
64'h3cc3c33cff00ff00,
64'hc33cc33cf0f0f0f0,
64'hc33cc33c0f0ff0f0,
64'h0ff00ff05a5a5a5a,
64'h5aa5a55a0ff00ff0,
64'hf00f0ff000ffff00,
64'hf0f0f0f03333cccc,
64'h6996699699996666,
64'h00000000ff00ff00,
64'h96696996f0f0f0f0,
64'hcc3333cca55aa55a,
64'hf00f0ff000ffff00,
64'hccccccccf00f0ff0,
64'h00000000cc3333cc,
64'h9966996633cc33cc,
64'h66666666aa5555aa,
64'h6969969666999966,
64'h66666666a55aa55a,
64'h000000003c3c3c3c,
64'hc33cc33c00ffff00,
64'h33cc33cc99996666,
64'h6969969669699696,
64'haa5555aa69699696,
64'h99669966cccccccc,
64'h33cc33cc66999966,
64'hcccccccc96696996,
64'h0ff00ff069966996,
64'hc3c33c3c5aa5a55a,
64'h3c3c3c3cc3c33c3c,
64'h00000000aaaaaaaa,
64'hcccccccc66999966,
64'h9669699696696996,
64'h6996699600ffff00,
64'h3333cccc00000000,
64'h0ff00ff05555aaaa,
64'h9966996633cc33cc,
64'ha55aa55a69699696,
64'h96969696c33cc33c,
64'h96969696f0f0f0f0,
64'h3cc3c33c3c3c3c3c,
64'h00ffff005555aaaa,
64'hc33cc33c5555aaaa,
64'hffff0000cc3333cc,
64'hcccccccc33cc33cc,
64'h96969696c3c33c3c,
64'h966969960f0ff0f0,
64'hffff000000000000,
64'h00000000cc3333cc,
64'hc33cc33c55aa55aa,
64'h5aa5a55a00ffff00,
64'hffff000000000000,
64'h0ff00ff0ff00ff00,
64'h5a5a5a5aaaaaaaaa,
64'h5555aaaa0f0ff0f0,
64'haa5555aa5555aaaa,
64'haa5555aa66999966,
64'hffff0000c33cc33c,
64'h3cc3c33c3333cccc,
64'hf0f0f0f0c3c33c3c,
64'h0ff00ff096969696,
64'haaaaaaaa3cc3c33c,
64'h00ffff000ff00ff0,
64'hcc3333cc69966996,
64'h0ff00ff03333cccc,
64'ha55aa55a55aa55aa,
64'hc3c33c3cc33cc33c,
64'hff00ff00a55aa55a,
64'h3333cccc96969696,
64'ha55aa55aff00ff00,
64'h5555aaaa5aa5a55a,
64'h99996666f0f0f0f0,
64'hccccccccffff0000,
64'hc3c33c3cf0f0f0f0,
64'h0000000066666666,
64'hf0f0f0f0cc3333cc,
64'h6969969669966996,
64'hf00f0ff03c3c3c3c,
64'hc3c33c3c55aa55aa,
64'hff00ff00c3c33c3c,
64'ha5a55a5a0f0ff0f0,
64'h55aa55aacc3333cc,
64'ha55aa55aff00ff00,
64'hffff000096696996,
64'h55aa55aa5555aaaa,
64'hc3c33c3c5aa5a55a,
64'h966969965555aaaa,
64'h00ffff0066666666,
64'haa5555aa5aa5a55a,
64'h5aa5a55a3c3c3c3c,
64'h9966996600000000,
64'h5aa5a55af0f0f0f0,
64'h0ff00ff066666666,
64'h33cc33cc5a5a5a5a,
64'h0000000033cc33cc,
64'h6699996600ffff00,
64'h99669966cc3333cc,
64'h33cc33cca5a55a5a,
64'h3cc3c33c00ffff00,
64'haaaaaaaa96696996,
64'hc3c33c3ca5a55a5a,
64'h00ffff0000000000,
64'h99996666ff00ff00,
64'h69699696c33cc33c,
64'hf0f0f0f03333cccc,
64'h55aa55aa3c3c3c3c,
64'h5555aaaaf00f0ff0,
64'h000000005aa5a55a,
64'hffff00005555aaaa,
64'hcc3333cc66666666,
64'ha5a55a5aa5a55a5a,
64'h3c3c3c3cff00ff00,
64'h9696969699996666,
64'hc33cc33c33cc33cc,
64'ha5a55a5a00000000,
64'h6996699666999966,
64'h33cc33cc66999966,
64'h0ff00ff03333cccc,
64'h96969696a55aa55a,
64'ha5a55a5a00000000,
64'hffff00003cc3c33c,
64'hc33cc33c5aa5a55a,
64'h5a5a5a5a69966996,
64'hc33cc33c0ff00ff0,
64'h6666666699996666,
64'hff00ff00cc3333cc,
64'hffff0000aa5555aa,
64'hffff0000c33cc33c,
64'h99669966cccccccc,
64'haa5555aa3333cccc,
64'h00ffff00c3c33c3c,
64'h6666666666666666,
64'hf00f0ff0ff00ff00,
64'hcc3333ccffff0000,
64'hcccccccc3c3c3c3c,
64'hc33cc33c3333cccc,
64'h9696969655aa55aa,
64'h96696996cccccccc,
64'h5a5a5a5a96696996,
64'ha5a55a5acc3333cc,
64'h33cc33cc3cc3c33c,
64'hf0f0f0f0cccccccc,
64'h5a5a5a5aff00ff00,
64'hffff00005555aaaa,
64'haaaaaaaaa5a55a5a,
64'h969696963c3c3c3c,
64'h0f0ff0f069966996,
64'h00ffff003c3c3c3c,
64'h6969969696696996,
64'h5aa5a55a69699696,
64'hc33cc33cf00f0ff0,
64'hffff00000f0ff0f0,
64'hcc3333cc66999966,
64'h3c3c3c3c5555aaaa,
64'h5aa5a55acc3333cc,
64'h3cc3c33c69699696,
64'h0f0ff0f0f0f0f0f0,
64'h33cc33ccc33cc33c,
64'h00ffff00cccccccc,
64'hffff000069966996,
64'h00000000c3c33c3c,
64'hc33cc33cf00f0ff0,
64'h33cc33cc33cc33cc,
64'h0ff00ff05a5a5a5a,
64'hf00f0ff00ff00ff0,
64'h00ffff0096969696,
64'hc33cc33c0ff00ff0,
64'h9966996633cc33cc,
64'h5a5a5a5a00ffff00,
64'h3c3c3c3ccccccccc,
64'hffff000096969696,
64'haaaaaaaaa5a55a5a,
64'h5aa5a55a66666666,
64'h5555aaaa33cc33cc,
64'h5a5a5a5ac33cc33c,
64'h9696969666666666,
64'hcccccccc3c3c3c3c,
64'h5a5a5a5a3cc3c33c,
64'h5aa5a55a55aa55aa,
64'hf0f0f0f03333cccc,
64'h9696969600ffff00,
64'h3c3c3c3c3c3c3c3c,
64'h69699696cc3333cc,
64'h3cc3c33c00000000,
64'h55aa55aaa55aa55a,
64'h5555aaaa66666666,
64'hc33cc33caa5555aa,
64'h5a5a5a5a3c3c3c3c,
64'h96969696c33cc33c,
64'h3cc3c33c3c3c3c3c,
64'hffff000000000000,
64'h5a5a5a5a00ffff00,
64'h33cc33cc5555aaaa,
64'h99996666f0f0f0f0,
64'ha55aa55a5a5a5a5a,
64'h996699665a5a5a5a,
64'h3333cccc5a5a5a5a,
64'h69699696ffff0000,
64'haa5555aa66666666,
64'h3333cccc99669966,
64'h00ffff00c33cc33c,
64'h96696996f0f0f0f0,
64'h6666666669966996,
64'h3333cccca5a55a5a,
64'h00ffff00aaaaaaaa,
64'h0ff00ff0f00f0ff0,
64'hff00ff005555aaaa,
64'h00ffff00ff00ff00,
64'h3c3c3c3cff00ff00,
64'h6666666699669966,
64'hc33cc33c00ffff00,
64'h3333ccccffff0000,
64'ha5a55a5a5a5a5a5a,
64'hf0f0f0f096969696,
64'h966969965555aaaa,
64'h0f0ff0f0ff00ff00,
64'h66666666cc3333cc,
64'h3333ccccffff0000,
64'h66999966aa5555aa,
64'h96696996a5a55a5a,
64'hffff0000a5a55a5a,
64'h969696963333cccc,
64'h6666666669699696,
64'h3c3c3c3c66999966,
64'h000000000ff00ff0,
64'h3c3c3c3cffff0000,
64'ha55aa55a96969696,
64'hf00f0ff069966996,
64'h6699996669966996,
64'hc33cc33c5a5a5a5a,
64'ha55aa55ac3c33c3c,
64'h5a5a5a5a96696996,
64'hf00f0ff096696996,
64'h3cc3c33ccc3333cc,
64'hffff0000a55aa55a,
64'h9669699666666666,
64'h5a5a5a5ac3c33c3c,
64'h9966996696696996,
64'h5a5a5a5a5555aaaa,
64'ha5a55a5aaaaaaaaa,
64'hcccccccccccccccc,
64'hffff0000a5a55a5a,
64'haaaaaaaac33cc33c,
64'h0ff00ff0a55aa55a,
64'hc33cc33cff00ff00,
64'hf00f0ff00ff00ff0,
64'h5555aaaacccccccc,
64'h5aa5a55a66666666,
64'h00000000a5a55a5a,
64'h5a5a5a5aa5a55a5a,
64'hc33cc33c0ff00ff0,
64'h3cc3c33c55aa55aa,
64'haaaaaaaaaaaaaaaa,
64'haaaaaaaa0f0ff0f0,
64'hf00f0ff099996666,
64'hcc3333ccffff0000,
64'haaaaaaaaaaaaaaaa,
64'haa5555aaffff0000,
64'h33cc33cccccccccc,
64'hccccccccff00ff00,
64'h9999666666666666,
64'h9999666669699696,
64'haaaaaaaa5aa5a55a,
64'h5aa5a55af0f0f0f0,
64'h55aa55aaa55aa55a,
64'h00ffff0069966996,
64'hccccccccf00f0ff0,
64'hffff0000aa5555aa,
64'ha5a55a5a3cc3c33c,
64'haa5555aaf0f0f0f0,
64'hcc3333cc99996666,
64'h0ff00ff0f00f0ff0,
64'h5555aaaacc3333cc,
64'hf0f0f0f0c33cc33c,
64'h66999966ffff0000,
64'hcccccccccc3333cc,
64'h9696969655aa55aa,
64'h5a5a5a5a00000000,
64'h0ff00ff055aa55aa,
64'haaaaaaaa3c3c3c3c,
64'hff00ff000f0ff0f0,
64'hc33cc33c96696996,
64'haa5555aa0ff00ff0,
64'ha55aa55a3333cccc,
64'h5555aaaa0ff00ff0,
64'h33cc33cc55aa55aa,
64'h99996666a5a55a5a,
64'hcc3333cc5555aaaa,
64'h000000003cc3c33c,
64'h9999666666666666,
64'h0ff00ff066999966,
64'h9669699666666666,
64'h5555aaaa96969696,
64'h99996666cc3333cc,
64'h66999966a55aa55a,
64'h6969969600000000,
64'hcc3333ccff00ff00,
64'haa5555aa3c3c3c3c,
64'h0f0ff0f033cc33cc,
64'h000000000f0ff0f0,
64'hc3c33c3cffff0000,
64'h69699696a5a55a5a,
64'h0f0ff0f099669966,
64'hf00f0ff05555aaaa,
64'h6666666696696996,
64'h0ff00ff099669966,
64'h5555aaaaaaaaaaaa,
64'h96969696ffff0000,
64'h69966996f00f0ff0,
64'h55aa55aaf0f0f0f0,
64'h3333cccca55aa55a,
64'hcccccccc00ffff00,
64'haaaaaaaa66999966,
64'h0000000066666666,
64'ha5a55a5a96969696,
64'h9966996633cc33cc,
64'ha55aa55a5555aaaa,
64'hc33cc33c3c3c3c3c,
64'hf00f0ff0a5a55a5a,
64'h33cc33cc00000000,
64'h96696996c3c33c3c,
64'h0f0ff0f069699696,
64'h00ffff005a5a5a5a,
64'hc33cc33c66999966,
64'h33cc33cc00000000,
64'haaaaaaaaf00f0ff0,
64'h5aa5a55a66999966,
64'h33cc33cc96696996,
64'hf00f0ff000ffff00,
64'h3c3c3c3c3c3c3c3c,
64'hffff0000a5a55a5a,
64'h0000000099996666,
64'haaaaaaaa5aa5a55a,
64'h69699696f0f0f0f0,
64'h3333ccccf0f0f0f0,
64'h5555aaaaa55aa55a,
64'h9696969696969696,
64'h00ffff00ffff0000,
64'ha5a55a5a00000000,
64'h5a5a5a5aa55aa55a,
64'hf00f0ff0f0f0f0f0,
64'hc33cc33c99996666,
64'h3cc3c33cf0f0f0f0,
64'h996699663cc3c33c,
64'h33cc33cca5a55a5a,
64'ha5a55a5a5aa5a55a,
64'hff00ff005a5a5a5a,
64'h33cc33ccffff0000,
64'h00000000cccccccc,
64'h6666666699669966,
64'hc33cc33ca55aa55a,
64'hff00ff003cc3c33c,
64'h5555aaaa0ff00ff0,
64'h699669963cc3c33c,
64'h6699996669966996,
64'h5aa5a55aaa5555aa,
64'h0000000055aa55aa,
64'ha5a55a5a69699696,
64'ha55aa55a66666666,
64'hcc3333cca5a55a5a,
64'h5aa5a55a69966996,
64'h55aa55aa55aa55aa,
64'ha5a55a5af00f0ff0,
64'hffff0000f0f0f0f0,
64'haaaaaaaa3cc3c33c,
64'haaaaaaaa0ff00ff0,
64'hf00f0ff0aa5555aa,
64'h0f0ff0f0a5a55a5a,
64'h00ffff0033cc33cc,
64'h00ffff0000ffff00,
64'h5555aaaac33cc33c,
64'h5aa5a55a00ffff00,
64'hc3c33c3c0f0ff0f0,
64'h33cc33ccffff0000,
64'h0ff00ff05a5a5a5a,
64'h00000000c33cc33c,
64'h6666666633cc33cc,
64'hcc3333cc96969696,
64'h666666660f0ff0f0,
64'h99669966f00f0ff0,
64'hc33cc33c3c3c3c3c,
64'hf0f0f0f00ff00ff0,
64'h33cc33ccf00f0ff0,
64'hcc3333cc99996666,
64'h55aa55aaf0f0f0f0,
64'hc33cc33c5555aaaa,
64'h0ff00ff0a55aa55a,
64'hc33cc33c0f0ff0f0,
64'h5aa5a55aaaaaaaaa,
64'h99996666cc3333cc,
64'hcccccccc3c3c3c3c,
64'h5aa5a55a3333cccc,
64'h33cc33cca55aa55a,
64'hc33cc33cf00f0ff0,
64'hf00f0ff00ff00ff0,
64'haaaaaaaa00000000,
64'h99669966ffff0000,
64'h0f0ff0f066666666,
64'h3c3c3c3c55aa55aa,
64'h6699996633cc33cc,
64'hc3c33c3c33cc33cc,
64'hf0f0f0f033cc33cc,
64'h6996699600000000,
64'h9999666696969696,
64'h5a5a5a5ac3c33c3c,
64'h5555aaaaf00f0ff0,
64'h96696996ff00ff00,
64'h969696963cc3c33c,
64'hf0f0f0f033cc33cc,
64'h5555aaaa66666666,
64'haa5555aa00ffff00,
64'hffff000066666666,
64'hffff00005555aaaa,
64'ha55aa55affff0000,
64'h3c3c3c3cc3c33c3c,
64'hf00f0ff0ffff0000,
64'hf0f0f0f0aaaaaaaa,
64'h9966996699669966,
64'h55aa55aac33cc33c,
64'h3cc3c33ccccccccc,
64'h55aa55aa5555aaaa,
64'h969696960f0ff0f0,
64'hf0f0f0f0aaaaaaaa,
64'h6969969699996666,
64'h9669699699669966,
64'haaaaaaaa99669966,
64'h699669965a5a5a5a,
64'h3c3c3c3c69966996,
64'h0ff00ff069699696,
64'h00000000aa5555aa,
64'h0ff00ff000000000,
64'hcc3333cc69966996,
64'h00ffff003cc3c33c,
64'h696996963cc3c33c,
64'h5aa5a55a33cc33cc,
64'hcc3333cc0ff00ff0,
64'h33cc33cc96696996,
64'h00ffff0096696996,
64'h5aa5a55aa5a55a5a,
64'haaaaaaaa66999966,
64'h966969963c3c3c3c,
64'h996699660ff00ff0,
64'hc3c33c3c96696996,
64'h33cc33cc66666666,
64'h33cc33cc66666666,
64'h5a5a5a5af0f0f0f0,
64'h0000000033cc33cc,
64'h666666665aa5a55a,
64'hff00ff0033cc33cc,
64'h5aa5a55affff0000,
64'h33cc33cc00ffff00,
64'h3c3c3c3cf0f0f0f0,
64'haa5555aa3c3c3c3c,
64'h5555aaaa33cc33cc,
64'h5555aaaa99669966,
64'h99669966aa5555aa,
64'h00ffff003333cccc,
64'h99996666cccccccc,
64'h69966996ff00ff00,
64'haaaaaaaa96969696,
64'hf00f0ff0aaaaaaaa,
64'hff00ff0066666666,
64'h5aa5a55a00000000,
64'haa5555aa5a5a5a5a,
64'h0f0ff0f0ffff0000,
64'h00ffff003c3c3c3c,
64'hccccccccc33cc33c,
64'h9999666666999966,
64'h5a5a5a5a55aa55aa,
64'h55aa55aacc3333cc,
64'h3333cccc3cc3c33c,
64'h3cc3c33c00ffff00,
64'h3cc3c33c99996666,
64'h666666665aa5a55a,
64'hf00f0ff055aa55aa,
64'haaaaaaaa3c3c3c3c,
64'h3cc3c33caa5555aa,
64'hcc3333cca5a55a5a,
64'haa5555aa5aa5a55a,
64'h0f0ff0f000000000,
64'hc33cc33ca5a55a5a,
64'hff00ff0099996666,
64'hf00f0ff000000000,
64'h966969963333cccc,
64'hcccccccc0ff00ff0,
64'hf00f0ff0ff00ff00,
64'hc3c33c3c96696996,
64'ha55aa55aaa5555aa,
64'h96969696f0f0f0f0,
64'h0ff00ff0aa5555aa,
64'h55aa55aa3333cccc,
64'h9999666633cc33cc,
64'h6969969666666666,
64'h5555aaaa5aa5a55a,
64'hff00ff0096969696,
64'hff00ff00c3c33c3c,
64'hcc3333cc96969696,
64'h99669966c33cc33c,
64'h699669960f0ff0f0,
64'h9999666666999966,
64'hcc3333cc00000000,
64'h96969696ffff0000,
64'h33cc33cc0ff00ff0,
64'h5555aaaa0f0ff0f0,
64'h69699696ff00ff00,
64'hf0f0f0f0aaaaaaaa,
64'haaaaaaaa99669966,
64'hf00f0ff069699696,
64'h3c3c3c3ccccccccc,
64'h33cc33cc96696996,
64'h55aa55aa69699696,
64'h96969696cccccccc,
64'h3333cccc00000000,
64'haa5555aaaa5555aa,
64'h3cc3c33c55aa55aa,
64'hf00f0ff0cc3333cc,
64'h00ffff00ffff0000,
64'h0f0ff0f069699696,
64'h5aa5a55a96969696,
64'hccccccccc33cc33c,
64'h996699660f0ff0f0,
64'hc3c33c3ccccccccc,
64'h3c3c3c3ca55aa55a,
64'h0ff00ff033cc33cc,
64'h96696996aaaaaaaa,
64'hf00f0ff00ff00ff0,
64'h9696969669966996,
64'h3cc3c33c99669966,
64'h96969696c3c33c3c,
64'h5a5a5a5aaaaaaaaa,
64'h9669699600ffff00,
64'hc33cc33c69699696,
64'h6996699696696996,
64'h0ff00ff05555aaaa,
64'ha55aa55aa55aa55a,
64'h00ffff0033cc33cc,
64'h9696969696969696,
64'h3333cccc66999966,
64'hc3c33c3c55aa55aa,
64'h00000000ff00ff00,
64'h99669966cc3333cc,
64'haa5555aac33cc33c,
64'haa5555aa00000000,
64'hc33cc33caaaaaaaa,
64'h5aa5a55acc3333cc,
64'h69699696ff00ff00,
64'h969696963c3c3c3c,
64'h6666666655aa55aa,
64'hc3c33c3cf00f0ff0,
64'h9999666699669966,
64'hf0f0f0f066999966,
64'h3c3c3c3c99669966,
64'hc33cc33c00000000,
64'h3c3c3c3c5a5a5a5a,
64'h5aa5a55ac3c33c3c,
64'h99669966cc3333cc,
64'haaaaaaaaf00f0ff0,
64'h96969696aa5555aa,
64'hc33cc33cf00f0ff0,
64'hf0f0f0f096696996,
64'h0f0ff0f03333cccc,
64'h33cc33cc99996666,
64'h69966996c33cc33c,
64'haaaaaaaa96969696,
64'h5aa5a55a33cc33cc,
64'h3333cccc96696996,
64'h0f0ff0f03333cccc,
64'hf0f0f0f000ffff00,
64'h3333cccc55aa55aa,
64'h3cc3c33cf00f0ff0,
64'h0f0ff0f0aa5555aa,
64'h696996963333cccc,
64'hf00f0ff099669966,
64'hff00ff00a5a55a5a,
64'h66666666ffff0000,
64'h3c3c3c3c5aa5a55a,
64'haa5555aaffff0000,
64'h00ffff0055aa55aa,
64'h69966996aaaaaaaa,
64'h0f0ff0f099669966,
64'h99669966f00f0ff0,
64'h3c3c3c3c0f0ff0f0,
64'h99669966c33cc33c,
64'hcc3333ccff00ff00,
64'h69699696aa5555aa,
64'h5aa5a55aa55aa55a,
64'h3cc3c33c00ffff00,
64'hc33cc33c00ffff00,
64'h5aa5a55a96969696,
64'hf0f0f0f055aa55aa,
64'hffff0000cccccccc,
64'haa5555aa66999966,
64'ha55aa55aff00ff00,
64'h5a5a5a5a66666666,
64'h3333cccc0f0ff0f0,
64'h66666666a55aa55a,
64'h00ffff00f0f0f0f0,
64'hcccccccc66999966,
64'hffff000000ffff00,
64'h5555aaaaaa5555aa,
64'hff00ff0000000000,
64'hcc3333cc00000000,
64'h5aa5a55a96969696,
64'h5aa5a55a3333cccc,
64'h0f0ff0f00f0ff0f0,
64'h00ffff000f0ff0f0,
64'hcccccccc0f0ff0f0,
64'h0f0ff0f000000000,
64'hc33cc33cc33cc33c,
64'hc3c33c3c0ff00ff0,
64'hf00f0ff0aa5555aa,
64'h000000005555aaaa,
64'h0f0ff0f0f00f0ff0,
64'h00ffff00a5a55a5a,
64'h969696963c3c3c3c,
64'h96969696ffff0000,
64'h0f0ff0f096969696,
64'hf0f0f0f0cccccccc,
64'haaaaaaaaaaaaaaaa,
64'h69699696a55aa55a,
64'h0ff00ff0aaaaaaaa,
64'hcccccccc66666666,
64'h33cc33ccc3c33c3c,
64'hff00ff00f00f0ff0,
64'h66666666f0f0f0f0,
64'haa5555aacccccccc,
64'h00ffff0055aa55aa,
64'h6666666666666666,
64'hffff00003c3c3c3c,
64'h0000000069699696,
64'h5a5a5a5ac3c33c3c,
64'h9669699633cc33cc,
64'haaaaaaaa3cc3c33c,
64'haa5555aac33cc33c,
64'h0000000099996666,
64'hccccccccaaaaaaaa,
64'ha55aa55a3cc3c33c,
64'h66666666f00f0ff0,
64'h969696965aa5a55a,
64'hcccccccca5a55a5a,
64'h0ff00ff000ffff00,
64'h0f0ff0f03cc3c33c,
64'h0f0ff0f096696996,
64'h55aa55aa99669966,
64'h3cc3c33c69699696,
64'haaaaaaaaa55aa55a,
64'hc3c33c3c00ffff00,
64'haa5555aa3cc3c33c,
64'h6996699696969696,
64'h5a5a5a5a3c3c3c3c,
64'h5555aaaaff00ff00,
64'h3c3c3c3c0f0ff0f0,
64'h5aa5a55acc3333cc,
64'hcccccccc5a5a5a5a,
64'h6699996600000000,
64'h969696965555aaaa,
64'h55aa55aa55aa55aa,
64'hffff00000ff00ff0,
64'h999966660f0ff0f0,
64'h00ffff00c3c33c3c,
64'h000000003333cccc,
64'h0f0ff0f05a5a5a5a,
64'h696996965a5a5a5a,
64'h3333ccccffff0000,
64'h66999966c33cc33c,
64'h5555aaaacccccccc,
64'hcc3333cc3c3c3c3c,
64'ha5a55a5a00000000,
64'h9669699633cc33cc,
64'haa5555aa00000000,
64'h69966996a55aa55a,
64'h00000000f00f0ff0,
64'hc3c33c3cc3c33c3c,
64'h0f0ff0f099996666,
64'hff00ff000f0ff0f0,
64'h3c3c3c3c5aa5a55a,
64'h3c3c3c3c5555aaaa,
64'h6666666696969696,
64'h6996699666999966,
64'h6969969699996666,
64'h696996960ff00ff0,
64'h669999663333cccc,
64'ha55aa55a99669966,
64'h6666666666999966,
64'h99669966aaaaaaaa,
64'hc3c33c3c33cc33cc,
64'hc3c33c3c96969696,
64'hc33cc33caaaaaaaa,
64'h00ffff00f0f0f0f0,
64'h5a5a5a5aaa5555aa,
64'h0f0ff0f0ffff0000,
64'h969696963cc3c33c,
64'hf0f0f0f099996666,
64'h3333cccc55aa55aa,
64'hc3c33c3c3333cccc,
64'hc33cc33c5a5a5a5a,
64'h99996666a5a55a5a,
64'ha55aa55a3c3c3c3c,
64'h99996666cc3333cc,
64'h9669699669966996,
64'haaaaaaaa0ff00ff0,
64'hffff000069966996,
64'h96696996f00f0ff0,
64'hc3c33c3cff00ff00,
64'hcccccccc69699696,
64'h00000000aaaaaaaa,
64'h5aa5a55a00000000,
64'ha55aa55aaa5555aa,
64'hcc3333ccff00ff00,
64'haa5555aa5555aaaa,
64'haaaaaaaacccccccc,
64'h0ff00ff0c3c33c3c,
64'ha55aa55ac33cc33c,
64'h3333cccc5a5a5a5a,
64'haa5555aa3cc3c33c,
64'h6666666669966996,
64'h996699665a5a5a5a,
64'haa5555aa00000000,
64'h0f0ff0f03333cccc,
64'h5555aaaa99996666,
64'haaaaaaaa0f0ff0f0,
64'h0ff00ff0aaaaaaaa,
64'h9669699669966996,
64'h3c3c3c3c69966996,
64'ha55aa55af00f0ff0,
64'h33cc33ccff00ff00,
64'h000000005a5a5a5a,
64'h69699696cc3333cc,
64'h0ff00ff00f0ff0f0,
64'h0f0ff0f0cccccccc,
64'h6699996600ffff00,
64'haaaaaaaa3cc3c33c,
64'h99996666c3c33c3c,
64'ha5a55a5a0ff00ff0,
64'h6699996666666666,
64'h66666666ffff0000,
64'h55aa55aa69966996,
64'hf0f0f0f096696996,
64'h0ff00ff066666666,
64'hcc3333cc66999966,
64'hff00ff000f0ff0f0,
64'h55aa55aac33cc33c,
64'h0f0ff0f0c3c33c3c,
64'ha5a55a5a99996666,
64'hf0f0f0f0ffff0000,
64'h3cc3c33c0f0ff0f0,
64'hf0f0f0f05aa5a55a,
64'hcc3333cc00000000,
64'h00ffff00cccccccc,
64'h0ff00ff00f0ff0f0,
64'h000000005555aaaa,
64'ha5a55a5a0ff00ff0,
64'haa5555aa3333cccc,
64'ha55aa55a00ffff00,
64'h0000000069699696,
64'h96969696c3c33c3c,
64'h6699996669699696,
64'h3c3c3c3c00000000,
64'h33cc33cc33cc33cc,
64'haaaaaaaa0ff00ff0,
64'h00000000a5a55a5a,
64'h99996666aa5555aa,
64'h9966996699996666,
64'ha55aa55aaa5555aa,
64'hcc3333cc96696996,
64'h969696965a5a5a5a,
64'h3cc3c33c96969696,
64'h669999665aa5a55a,
64'h00ffff00c33cc33c,
64'h999966660f0ff0f0,
64'h0ff00ff03cc3c33c,
64'hc33cc33c5a5a5a5a,
64'h969696965555aaaa,
64'h6969969699996666,
64'h0000000000ffff00,
64'h9669699699996666,
64'h000000005a5a5a5a,
64'h0ff00ff069699696,
64'hff00ff0033cc33cc,
64'h0f0ff0f0aaaaaaaa,
64'h55aa55aa66999966,
64'hffff0000aaaaaaaa,
64'hf0f0f0f099996666,
64'h5a5a5a5acccccccc,
64'hf0f0f0f0c3c33c3c,
64'hf00f0ff000ffff00,
64'h0ff00ff055aa55aa,
64'h55aa55aa5aa5a55a,
64'h55aa55aaffff0000,
64'hc33cc33c3333cccc,
64'hcc3333cc66999966,
64'h99669966ffff0000,
64'h969696965555aaaa,
64'h9999666669966996,
64'h3cc3c33c3333cccc,
64'h0ff00ff0f0f0f0f0,
64'h3333ccccc3c33c3c,
64'h33cc33cc5555aaaa,
64'ha5a55a5a3c3c3c3c,
64'h5555aaaaff00ff00,
64'haaaaaaaa66999966,
64'h3333ccccff00ff00,
64'h3333ccccc3c33c3c,
64'h0ff00ff05555aaaa,
64'h33cc33cc99996666,
64'hcc3333ccaaaaaaaa,
64'h00ffff0000000000,
64'hc33cc33cc33cc33c,
64'h99669966f0f0f0f0,
64'h9966996655aa55aa,
64'hf0f0f0f055aa55aa,
64'hc33cc33c55aa55aa,
64'hccccccccaaaaaaaa,
64'ha5a55a5af00f0ff0,
64'h5555aaaa00ffff00,
64'h969696963333cccc,
64'h3cc3c33c66666666,
64'h99996666aa5555aa,
64'haaaaaaaa99669966,
64'h33cc33cca55aa55a,
64'hcc3333cc00000000,
64'h5aa5a55a69966996,
64'h0ff00ff0f0f0f0f0,
64'h00ffff00cccccccc,
64'ha5a55a5acc3333cc,
64'ha55aa55acccccccc,
64'h699669963c3c3c3c,
64'hff00ff000ff00ff0,
64'h33cc33ccaa5555aa,
64'haa5555aa55aa55aa,
64'h00ffff00f0f0f0f0,
64'h969696963333cccc,
64'h0ff00ff03c3c3c3c,
64'h3cc3c33c0ff00ff0,
64'h3cc3c33cc33cc33c,
64'h0ff00ff0a55aa55a,
64'h96696996a5a55a5a,
64'hc33cc33cf00f0ff0,
64'h999966665aa5a55a,
64'haaaaaaaa3c3c3c3c,
64'h3cc3c33c66666666,
64'h66666666f00f0ff0,
64'h0f0ff0f0aa5555aa,
64'h3c3c3c3c66999966,
64'h5aa5a55a99669966,
64'haaaaaaaa5555aaaa,
64'h55aa55aa5aa5a55a,
64'ha55aa55a96696996,
64'haaaaaaaa69699696,
64'haaaaaaaac33cc33c,
64'hf00f0ff066999966,
64'ha55aa55affff0000,
64'h3c3c3c3c5aa5a55a,
64'h5a5a5a5a69966996,
64'h669999660ff00ff0,
64'haa5555aaffff0000,
64'h99669966ff00ff00,
64'haaaaaaaaa5a55a5a,
64'h9696969699669966,
64'hc3c33c3caaaaaaaa,
64'h69966996ffff0000,
64'h3333ccccc3c33c3c,
64'h00000000cc3333cc,
64'h9696969600ffff00,
64'h5555aaaac3c33c3c,
64'haaaaaaaa3333cccc,
64'hff00ff0069966996,
64'h69966996cc3333cc,
64'h5a5a5a5aa55aa55a,
64'h69699696f0f0f0f0,
64'h66666666a55aa55a,
64'ha5a55a5a96969696,
64'h9966996669966996,
64'h9669699600ffff00,
64'h99996666ffff0000,
64'h96696996f0f0f0f0,
64'h000000005aa5a55a,
64'h0ff00ff05aa5a55a,
64'h55aa55aa00ffff00,
64'h5555aaaa99996666,
64'h0ff00ff0aa5555aa,
64'h0ff00ff000ffff00,
64'h3c3c3c3c5555aaaa,
64'h3cc3c33c3cc3c33c,
64'hc33cc33cff00ff00,
64'h69966996a55aa55a,
64'h6969969666666666,
64'h6699996669966996,
64'h3c3c3c3c3c3c3c3c,
64'hc3c33c3caaaaaaaa,
64'h0ff00ff096696996,
64'ha55aa55aff00ff00,
64'h5aa5a55a0f0ff0f0,
64'hffff000069966996,
64'h996699663333cccc,
64'hff00ff00a55aa55a,
64'h6996699669699696,
64'hff00ff0000ffff00,
64'hf0f0f0f069966996,
64'ha55aa55a33cc33cc,
64'h5aa5a55a69699696,
64'h3c3c3c3c96696996,
64'h6699996669966996,
64'h3c3c3c3cf0f0f0f0,
64'h966969965555aaaa,
64'h6666666655aa55aa,
64'h00000000cc3333cc,
64'h96696996ffff0000,
64'ha55aa55aaa5555aa,
64'h5a5a5a5a33cc33cc,
64'h00000000c3c33c3c,
64'hcc3333cc3333cccc,
64'h6699996699669966,
64'h0f0ff0f055aa55aa,
64'h999966660f0ff0f0,
64'h66666666a55aa55a,
64'h00ffff00cccccccc,
64'hcc3333ccff00ff00,
64'hf0f0f0f0a5a55a5a,
64'h999966665555aaaa,
64'h96969696c33cc33c,
64'hc3c33c3c69966996,
64'h3333cccc5aa5a55a,
64'h55aa55aa66666666,
64'h6666666699669966,
64'h666666665555aaaa,
64'h00ffff003cc3c33c,
64'h3cc3c33cff00ff00,
64'ha55aa55a66666666,
64'hcc3333ccffff0000,
64'h0f0ff0f0a55aa55a,
64'h000000003c3c3c3c,
64'hc33cc33cc33cc33c,
64'haa5555aa5aa5a55a,
64'hff00ff0069966996,
64'h696996963333cccc,
64'h6666666699996666,
64'h3c3c3c3ccccccccc,
64'h9966996666666666,
64'h6969969669699696,
64'h969696965aa5a55a,
64'h3333cccc99669966,
64'hff00ff00f0f0f0f0,
64'h00ffff0099996666,
64'h0f0ff0f0c3c33c3c,
64'h5555aaaa5555aaaa,
64'h3333cccc66999966,
64'hff00ff00f00f0ff0,
64'h9966996696696996,
64'h55aa55aaf0f0f0f0,
64'hf00f0ff0aaaaaaaa,
64'h55aa55aaa55aa55a,
64'h0f0ff0f0ff00ff00,
64'h5555aaaaaaaaaaaa,
64'haa5555aa3cc3c33c,
64'h000000000ff00ff0,
64'h33cc33cc66666666,
64'h9999666666999966,
64'h66999966ffff0000,
64'h00000000ff00ff00,
64'hc33cc33c66666666,
64'hc3c33c3c00ffff00,
64'ha55aa55a66999966,
64'h0f0ff0f03333cccc,
64'hcccccccc66666666,
64'h000000005aa5a55a,
64'h3c3c3c3ccccccccc,
64'h69699696cccccccc,
64'hcc3333cccccccccc,
64'h0f0ff0f0a55aa55a,
64'h69966996f0f0f0f0,
64'hf00f0ff05a5a5a5a,
64'h6969969696696996,
64'h5555aaaa96969696,
64'h96969696aaaaaaaa,
64'haa5555aa0f0ff0f0,
64'hf00f0ff00ff00ff0,
64'hc33cc33c0ff00ff0,
64'hc33cc33c0f0ff0f0,
64'haaaaaaaa0ff00ff0,
64'h3cc3c33c5555aaaa,
64'haaaaaaaaf0f0f0f0,
64'h00ffff0066999966,
64'hffff00000ff00ff0,
64'hff00ff00ffff0000,
64'h9999666699996666,
64'h00000000aaaaaaaa,
64'h55aa55aa99996666,
64'h33cc33cc96696996,
64'hff00ff0000000000,
64'h00ffff00cc3333cc,
64'haa5555aa99996666,
64'h3333cccc5a5a5a5a,
64'h3333ccccf00f0ff0,
64'hf00f0ff0f0f0f0f0,
64'h0f0ff0f0c3c33c3c,
64'h6969969669699696,
64'hc33cc33caa5555aa,
64'h3c3c3c3cc3c33c3c,
64'h5aa5a55a99996666,
64'haa5555aa5a5a5a5a,
64'hf0f0f0f0a55aa55a,
64'ha5a55a5a3333cccc,
64'h33cc33cc3333cccc,
64'h666666665a5a5a5a,
64'h66666666ffff0000,
64'hf0f0f0f099996666,
64'h5a5a5a5a66999966,
64'haa5555aa69966996,
64'h0f0ff0f0c33cc33c,
64'h0f0ff0f0ff00ff00,
64'h5555aaaa0ff00ff0,
64'h5aa5a55a55aa55aa,
64'hc3c33c3c00ffff00,
64'hc3c33c3cffff0000,
64'hff00ff0096969696,
64'hf00f0ff0aa5555aa,
64'hf0f0f0f0ff00ff00,
64'h33cc33ccffff0000,
64'h666666660ff00ff0,
64'h6996699666999966,
64'hf00f0ff000ffff00,
64'h9696969655aa55aa,
64'h6666666696969696,
64'h0f0ff0f096696996,
64'h0f0ff0f00f0ff0f0,
64'h6699996699669966,
64'haa5555aaa55aa55a,
64'hffff00003cc3c33c,
64'h9966996669966996,
64'h669999665555aaaa,
64'h3cc3c33c96969696,
64'hffff0000f0f0f0f0,
64'h0f0ff0f0ff00ff00,
64'h3333cccc0ff00ff0,
64'h5555aaaacccccccc,
64'h699669963333cccc,
64'h00ffff003c3c3c3c,
64'hf00f0ff03c3c3c3c,
64'h5aa5a55a66666666,
64'haa5555aaf00f0ff0,
64'h3cc3c33c99669966,
64'h5aa5a55a0f0ff0f0,
64'h3c3c3c3ccc3333cc,
64'h66666666a55aa55a,
64'hf00f0ff0f00f0ff0,
64'h96969696aaaaaaaa,
64'hff00ff00aaaaaaaa,
64'ha55aa55a96696996,
64'hcc3333ccc33cc33c,
64'h6666666666999966,
64'h3333cccccc3333cc,
64'hcc3333cc66999966,
64'hcccccccc5aa5a55a,
64'hcccccccc00000000,
64'h00ffff0055aa55aa,
64'h6699996600000000,
64'h0ff00ff0c33cc33c,
64'h33cc33cc5a5a5a5a,
64'hc3c33c3c55aa55aa,
64'h9999666666999966,
64'h6969969669699696,
64'hcccccccc5555aaaa,
64'hc33cc33c5a5a5a5a,
64'ha55aa55a66666666,
64'ha55aa55a3333cccc,
64'haaaaaaaaff00ff00,
64'h6666666669699696,
64'h3cc3c33caaaaaaaa,
64'haa5555aac3c33c3c,
64'h0f0ff0f03333cccc,
64'h0f0ff0f066999966,
64'hc33cc33cf0f0f0f0,
64'h96969696c3c33c3c,
64'h696996965555aaaa,
64'hc33cc33c99996666,
64'haaaaaaaa5a5a5a5a,
64'h00ffff005555aaaa,
64'h3333ccccf00f0ff0,
64'h696996965555aaaa,
64'haaaaaaaa69699696,
64'hf0f0f0f096696996,
64'hff00ff0099669966,
64'ha55aa55ac33cc33c,
64'h00ffff005aa5a55a,
64'h669999665555aaaa,
64'h6666666633cc33cc,
64'h3333cccc5aa5a55a,
64'h0f0ff0f0a5a55a5a,
64'h3333cccc3cc3c33c,
64'h33cc33ccc33cc33c,
64'h55aa55aaaaaaaaaa,
64'h699669963c3c3c3c,
64'h5aa5a55af00f0ff0,
64'hc33cc33c00000000,
64'h3333cccca5a55a5a,
64'hf00f0ff069699696,
64'h0ff00ff03cc3c33c,
64'h3c3c3c3c00ffff00,
64'h69699696f0f0f0f0,
64'hf00f0ff069699696,
64'h0f0ff0f0f0f0f0f0,
64'h69966996c33cc33c,
64'h0f0ff0f066666666,
64'h0f0ff0f0cc3333cc,
64'h3c3c3c3c3333cccc,
64'h00ffff0033cc33cc,
64'h0f0ff0f05aa5a55a,
64'h5aa5a55a00ffff00,
64'hffff00000ff00ff0,
64'hc3c33c3ccccccccc,
64'hf0f0f0f0ffff0000,
64'hc3c33c3c55aa55aa,
64'h9999666666999966,
64'hc33cc33c5555aaaa,
64'ha5a55a5aaa5555aa,
64'h3c3c3c3c69699696,
64'hc33cc33cc33cc33c,
64'h5555aaaa33cc33cc,
64'h5555aaaa3cc3c33c,
64'h6996699699996666,
64'h3cc3c33c33cc33cc,
64'h000000005a5a5a5a,
64'hc3c33c3ca5a55a5a,
64'h99669966c33cc33c,
64'h3cc3c33c0ff00ff0,
64'h55aa55aa66999966,
64'h00ffff0096969696,
64'h0f0ff0f000000000,
64'h33cc33cccc3333cc,
64'h3cc3c33ccc3333cc,
64'ha55aa55a00000000,
64'h9966996696969696,
64'h3c3c3c3c66999966,
64'hf00f0ff0ff00ff00,
64'ha5a55a5a96969696,
64'ha55aa55a00000000,
64'h3c3c3c3c3c3c3c3c,
64'h3c3c3c3cc33cc33c,
64'h66999966a5a55a5a,
64'h0ff00ff03c3c3c3c,
64'h55aa55aa55aa55aa,
64'h6666666633cc33cc,
64'h0ff00ff0f00f0ff0,
64'h9669699696696996,
64'h3333cccc3c3c3c3c,
64'hffff000066666666,
64'h996699663333cccc,
64'hf0f0f0f03333cccc,
64'h55aa55aaa55aa55a,
64'h6699996666999966,
64'h666666665555aaaa,
64'haaaaaaaa55aa55aa,
64'hc33cc33c96969696,
64'h696996960ff00ff0,
64'hffff000033cc33cc,
64'h5a5a5a5a0ff00ff0,
64'haaaaaaaaaa5555aa,
64'h3c3c3c3c96969696,
64'h5a5a5a5a33cc33cc,
64'hc33cc33cc3c33c3c,
64'hc33cc33cf00f0ff0,
64'haa5555aa55aa55aa,
64'hc3c33c3c00000000,
64'h3c3c3c3cc3c33c3c,
64'h3333ccccff00ff00,
64'h6699996696969696,
64'haaaaaaaaa55aa55a,
64'hc33cc33c66666666,
64'h3cc3c33cf00f0ff0,
64'h69699696a55aa55a,
64'h5aa5a55a0f0ff0f0,
64'h99669966aaaaaaaa,
64'hf0f0f0f0a5a55a5a,
64'h66999966ff00ff00,
64'hffff000096969696,
64'h99996666aaaaaaaa,
64'h33cc33cc66999966,
64'haa5555aaa5a55a5a,
64'h3c3c3c3c99669966,
64'h66999966aaaaaaaa,
64'h3cc3c33c3cc3c33c,
64'h99996666c3c33c3c,
64'h6996699666999966,
64'h96696996f0f0f0f0,
64'h33cc33cc0f0ff0f0,
64'h0ff00ff03c3c3c3c,
64'h5a5a5a5a66666666,
64'h00ffff0000000000,
64'h666666663333cccc,
64'h66666666cccccccc,
64'h66666666aaaaaaaa,
64'h9696969699996666,
64'hc33cc33c5a5a5a5a,
64'hf00f0ff0a55aa55a,
64'h6699996696696996,
64'h9999666696969696,
64'hcc3333cc0f0ff0f0,
64'h00ffff005a5a5a5a,
64'h00ffff00ff00ff00,
64'hff00ff00a55aa55a,
64'haa5555aaaa5555aa,
64'h9696969655aa55aa,
64'h5a5a5a5af0f0f0f0,
64'ha55aa55affff0000,
64'h9669699696969696,
64'hff00ff0066999966,
64'h66999966a5a55a5a,
64'h33cc33cccc3333cc,
64'h999966663cc3c33c,
64'h000000003c3c3c3c,
64'h33cc33cc5a5a5a5a,
64'h5aa5a55a00000000,
64'h3cc3c33c99996666,
64'h00000000a5a55a5a,
64'hcccccccc66999966,
64'h699669960f0ff0f0,
64'hc33cc33c96969696,
64'h5aa5a55a00000000,
64'h6996699666666666,
64'hf0f0f0f0cc3333cc,
64'h99996666aa5555aa,
64'h6666666666999966,
64'hf00f0ff0ff00ff00,
64'h66999966f0f0f0f0,
64'h00000000ff00ff00,
64'h96969696c33cc33c,
64'h0f0ff0f0ff00ff00,
64'hc3c33c3c3cc3c33c,
64'ha55aa55a66999966,
64'h5aa5a55a5aa5a55a,
64'hcccccccccccccccc,
64'hc3c33c3c96696996,
64'h669999663c3c3c3c,
64'h0ff00ff0f0f0f0f0,
64'hccccccccc3c33c3c,
64'hc3c33c3cf0f0f0f0,
64'h5aa5a55a0f0ff0f0,
64'h9999666633cc33cc,
64'hcc3333cc96969696,
64'h55aa55aac33cc33c,
64'h55aa55aa3333cccc,
64'h669999663c3c3c3c,
64'h969696963333cccc,
64'hf0f0f0f0aa5555aa,
64'ha5a55a5a3cc3c33c,
64'hf00f0ff0c3c33c3c,
64'hc3c33c3c5a5a5a5a,
64'h0ff00ff00f0ff0f0,
64'h3c3c3c3c66999966,
64'hcccccccccccccccc,
64'hc3c33c3ccc3333cc,
64'hccccccccffff0000,
64'h3333ccccc3c33c3c,
64'ha55aa55af0f0f0f0,
64'h3cc3c33c69966996,
64'h5a5a5a5a0f0ff0f0,
64'h5555aaaa99996666,
64'h6969969655aa55aa,
64'haa5555aaf00f0ff0,
64'h69966996a55aa55a,
64'hc3c33c3caaaaaaaa,
64'h0ff00ff055aa55aa,
64'hc33cc33cffff0000,
64'h5aa5a55a66666666,
64'hf00f0ff0a55aa55a,
64'h55aa55aa55aa55aa,
64'h3cc3c33c00ffff00,
64'hc33cc33c55aa55aa,
64'h669999663c3c3c3c,
64'hff00ff00f0f0f0f0,
64'h969696965555aaaa,
64'hf0f0f0f0c33cc33c,
64'h0ff00ff066666666,
64'hff00ff000ff00ff0,
64'h3cc3c33c5a5a5a5a,
64'ha55aa55a69699696,
64'ha55aa55a55aa55aa,
64'h666666660ff00ff0,
64'h6969969666666666,
64'h0f0ff0f096969696,
64'h55aa55aa99669966,
64'h96696996cccccccc,
64'h55aa55aaaa5555aa,
64'h9669699666666666,
64'h5aa5a55a69966996,
64'ha55aa55a96696996,
64'h0000000069699696,
64'h5a5a5a5af00f0ff0,
64'h33cc33cccc3333cc,
64'ha5a55a5a66666666,
64'hf00f0ff0a5a55a5a,
64'hcc3333cccc3333cc,
64'haaaaaaaa99669966,
64'h33cc33cc5aa5a55a,
64'haaaaaaaa5aa5a55a,
64'ha5a55a5acccccccc,
64'h3c3c3c3c0ff00ff0,
64'h33cc33cc00ffff00,
64'h96696996aaaaaaaa,
64'h6996699633cc33cc,
64'h9669699669966996,
64'h699669965aa5a55a,
64'h996699665555aaaa,
64'hc33cc33c55aa55aa,
64'ha5a55a5ac33cc33c,
64'h6666666655aa55aa,
64'h00000000f00f0ff0,
64'h0f0ff0f03c3c3c3c,
64'h969696960f0ff0f0,
64'h5555aaaa5a5a5a5a,
64'h5a5a5a5aa5a55a5a,
64'h99669966cc3333cc,
64'h996699665555aaaa,
64'h69966996aa5555aa,
64'hf00f0ff0f0f0f0f0,
64'ha55aa55a00000000,
64'hf0f0f0f099996666,
64'h69966996c3c33c3c,
64'haa5555aa66666666,
64'h9669699699996666,
64'h9669699669966996,
64'h5a5a5a5a5aa5a55a,
64'hcc3333cc0f0ff0f0,
64'ha5a55a5af00f0ff0,
64'h6969969696969696,
64'h3333cccca5a55a5a,
64'h0f0ff0f033cc33cc,
64'h9999666633cc33cc,
64'hcc3333cc5aa5a55a,
64'ha55aa55a00ffff00,
64'hc3c33c3cc3c33c3c,
64'ha55aa55a69966996,
64'hc33cc33c00000000,
64'haa5555aa0f0ff0f0,
64'hf0f0f0f0a5a55a5a,
64'h3c3c3c3caaaaaaaa,
64'h00000000c33cc33c,
64'h5555aaaac3c33c3c,
64'hffff00005555aaaa,
64'h69699696c33cc33c,
64'h6969969600000000,
64'hc3c33c3c0ff00ff0,
64'h00ffff00f00f0ff0,
64'hf00f0ff033cc33cc,
64'h66999966a55aa55a,
64'hf00f0ff03333cccc,
64'h55aa55aa0f0ff0f0,
64'hcccccccc00ffff00,
64'h6996699696696996,
64'h00ffff00a55aa55a,
64'ha5a55a5a3c3c3c3c,
64'ha55aa55af0f0f0f0,
64'hf00f0ff05a5a5a5a,
64'h3333cccc66999966,
64'hc33cc33cc3c33c3c,
64'haaaaaaaa66666666,
64'h3333cccc99996666,
64'hf0f0f0f0c33cc33c,
64'h9966996600ffff00,
64'h55aa55aa0f0ff0f0,
64'h5aa5a55a00ffff00,
64'h996699663333cccc,
64'h55aa55aa69966996,
64'hf00f0ff00f0ff0f0,
64'h999966660ff00ff0,
64'h3c3c3c3caa5555aa,
64'ha55aa55a99996666,
64'h0ff00ff000000000,
64'h33cc33cc0ff00ff0,
64'h33cc33cc5555aaaa,
64'h00000000c33cc33c,
64'haa5555aacc3333cc,
64'hcc3333cc3c3c3c3c,
64'h9696969600ffff00,
64'h00ffff0066999966,
64'h33cc33ccff00ff00,
64'h3333cccc66666666,
64'haa5555aa33cc33cc,
64'hf0f0f0f05555aaaa,
64'hc33cc33cc33cc33c,
64'h0ff00ff0cccccccc,
64'hffff0000c3c33c3c,
64'hff00ff0099669966,
64'hf0f0f0f069699696,
64'h96696996cccccccc,
64'hcc3333ccf00f0ff0,
64'h55aa55aaa55aa55a,
64'h0ff00ff069699696,
64'h6666666655aa55aa,
64'h66666666ff00ff00,
64'h69699696a55aa55a,
64'h966969963c3c3c3c,
64'h55aa55aa00000000,
64'ha5a55a5af0f0f0f0,
64'h666666665a5a5a5a,
64'hf0f0f0f0cccccccc,
64'h669999663c3c3c3c,
64'h3c3c3c3c99669966,
64'h0f0ff0f0cc3333cc,
64'hf00f0ff03cc3c33c,
64'h9696969669966996,
64'h33cc33ccff00ff00,
64'h0ff00ff099669966,
64'hffff0000ffff0000,
64'hffff0000cc3333cc,
64'hf0f0f0f03333cccc,
64'ha5a55a5a99996666,
64'h66666666ff00ff00,
64'ha55aa55a00000000,
64'h3333cccc69966996,
64'hffff0000c3c33c3c,
64'h9696969699669966,
64'h33cc33cca5a55a5a,
64'h999966665aa5a55a,
64'h96969696a55aa55a,
64'hc3c33c3c33cc33cc,
64'ha55aa55a00000000,
64'h5555aaaa3c3c3c3c,
64'hff00ff0099669966,
64'h6996699669699696,
64'h3333cccc55aa55aa,
64'h55aa55aa69966996,
64'h33cc33cc00000000,
64'h5aa5a55a3c3c3c3c,
64'h5aa5a55a0f0ff0f0,
64'ha55aa55a99996666,
64'ha55aa55a69699696,
64'hffff00005555aaaa,
64'h33cc33ccff00ff00,
64'h96696996ffff0000,
64'h5555aaaaf00f0ff0,
64'h99996666ffff0000,
64'h5aa5a55af00f0ff0,
64'h3cc3c33c69699696,
64'hc33cc33c66999966,
64'hffff00005a5a5a5a,
64'h55aa55aa3cc3c33c,
64'ha55aa55aa55aa55a,
64'hccccccccff00ff00,
64'hffff00000ff00ff0,
64'h9696969655aa55aa,
64'h96969696ff00ff00,
64'h5aa5a55aa5a55a5a,
64'h33cc33ccc33cc33c,
64'haa5555aaf00f0ff0,
64'hf0f0f0f0f0f0f0f0,
64'h5aa5a55aa55aa55a,
64'h5555aaaaf0f0f0f0,
64'h6969969699996666,
64'h0ff00ff05aa5a55a,
64'h00ffff00a55aa55a,
64'h0000000099669966,
64'h00ffff00ff00ff00,
64'h0ff00ff069699696,
64'h3cc3c33c5a5a5a5a,
64'ha5a55a5a0f0ff0f0,
64'h69699696aaaaaaaa,
64'h0ff00ff0a55aa55a,
64'hcccccccc55aa55aa,
64'h5a5a5a5a3cc3c33c,
64'h33cc33ccff00ff00,
64'h3c3c3c3c96969696,
64'h5aa5a55a99996666,
64'hc33cc33c00ffff00,
64'h0000000066999966,
64'ha55aa55acccccccc,
64'h0ff00ff03333cccc,
64'h3c3c3c3c00000000,
64'h9966996696969696,
64'hcccccccccc3333cc,
64'ha5a55a5a3333cccc,
64'h96969696ffff0000,
64'h6996699666666666,
64'hc3c33c3c0ff00ff0,
64'h5555aaaaff00ff00,
64'hc33cc33ccccccccc,
64'hff00ff005aa5a55a,
64'h00ffff003c3c3c3c,
64'hffff000000ffff00,
64'hf00f0ff033cc33cc,
64'h66999966c33cc33c,
64'hcc3333cc99996666,
64'h3c3c3c3c00ffff00,
64'hc33cc33c3c3c3c3c,
64'h55aa55aac33cc33c,
64'h99996666c3c33c3c,
64'h3cc3c33cf0f0f0f0,
64'h999966663333cccc,
64'h3cc3c33c96969696,
64'h669999663cc3c33c,
64'h669999663cc3c33c,
64'h0000000069966996,
64'h33cc33ccaa5555aa,
64'h0f0ff0f0a5a55a5a,
64'h33cc33cc96969696,
64'haa5555aa33cc33cc,
64'ha5a55a5aa5a55a5a,
64'h6666666669699696,
64'h0f0ff0f0cc3333cc,
64'hcccccccc66999966,
64'h33cc33cc5a5a5a5a,
64'ha55aa55a00ffff00,
64'h0f0ff0f0ffff0000,
64'h3cc3c33c66666666,
64'h966969960f0ff0f0,
64'h3cc3c33c3cc3c33c,
64'h96696996cc3333cc,
64'hc3c33c3c66666666,
64'hf00f0ff099996666,
64'h33cc33ccf00f0ff0,
64'h969696963333cccc,
64'h0000000000ffff00,
64'hff00ff00a55aa55a,
64'h69966996ff00ff00,
64'hcccccccc99669966,
64'h9966996633cc33cc,
64'hc3c33c3ca5a55a5a,
64'hc3c33c3c66666666,
64'h3cc3c33c99996666,
64'h00ffff0055aa55aa,
64'h6699996600000000,
64'hff00ff003c3c3c3c,
64'h3cc3c33ca55aa55a,
64'h3333cccc96969696,
64'h966969963c3c3c3c,
64'h9669699696696996,
64'h99669966cc3333cc,
64'h0f0ff0f055aa55aa,
64'h99669966aa5555aa,
64'h6996699669966996,
64'h5a5a5a5a33cc33cc,
64'h55aa55aaa5a55a5a,
64'h969696960f0ff0f0,
64'ha5a55a5acc3333cc,
64'h669999665555aaaa,
64'h0ff00ff0a55aa55a,
64'h6699996696696996,
64'hf00f0ff000000000,
64'h3333ccccff00ff00,
64'h55aa55aa99669966,
64'h0ff00ff066666666,
64'h00000000f00f0ff0,
64'hcccccccc0ff00ff0,
64'haaaaaaaa66666666,
64'h699669965aa5a55a,
64'h6996699600000000,
64'ha55aa55a00ffff00,
64'h5555aaaa00ffff00,
64'haa5555aaa5a55a5a,
64'h69699696cc3333cc,
64'haa5555aaf0f0f0f0,
64'h9999666655aa55aa,
64'hf0f0f0f05555aaaa,
64'h3cc3c33c96696996,
64'hffff000066999966,
64'h996699660ff00ff0,
64'h66999966ff00ff00,
64'h00ffff0033cc33cc,
64'h5a5a5a5ac3c33c3c,
64'h5aa5a55aa55aa55a,
64'hcccccccc96969696,
64'hf0f0f0f03c3c3c3c,
64'h55aa55aa5aa5a55a,
64'hc3c33c3cffff0000,
64'h3333cccc55aa55aa,
64'hcc3333cc5555aaaa,
64'h696996965a5a5a5a,
64'h3333cccc96696996,
64'h00ffff00ff00ff00,
64'h96969696aa5555aa,
64'ha55aa55a3333cccc,
64'hcc3333cc96969696,
64'h00ffff00aaaaaaaa,
64'h0f0ff0f000ffff00,
64'h0f0ff0f0cccccccc,
64'h000000005aa5a55a,
64'h3333cccc0f0ff0f0,
64'ha5a55a5aa55aa55a,
64'h69966996ffff0000,
64'hffff000069699696,
64'ha5a55a5a5555aaaa,
64'hf0f0f0f03c3c3c3c,
64'h999966660f0ff0f0,
64'h55aa55aacccccccc,
64'hf00f0ff05aa5a55a,
64'h00ffff00f0f0f0f0,
64'h000000000ff00ff0,
64'h5555aaaa69699696,
64'hff00ff00c33cc33c,
64'h3cc3c33c5a5a5a5a,
64'ha5a55a5a00ffff00,
64'h9999666666999966,
64'h00ffff00c33cc33c,
64'h3c3c3c3c99996666,
64'h3c3c3c3cffff0000,
64'hc33cc33ccc3333cc,
64'h966969960ff00ff0,
64'h9999666600000000,
64'h33cc33ccff00ff00,
64'h9696969633cc33cc,
64'hff00ff00f0f0f0f0,
64'hc3c33c3c0ff00ff0,
64'ha55aa55ac3c33c3c,
64'hff00ff000f0ff0f0,
64'haa5555aa5aa5a55a,
64'h6996699696696996,
64'h0f0ff0f0ffff0000,
64'h00ffff00c3c33c3c,
64'h0000000000000000,
64'haaaaaaaaa5a55a5a,
64'h55aa55aa5a5a5a5a,
64'h33cc33cc96969696,
64'h969696965555aaaa,
64'hcc3333cc00000000,
64'hf0f0f0f03cc3c33c,
64'haaaaaaaa0ff00ff0,
64'h6996699669699696,
64'h0f0ff0f033cc33cc,
64'h3c3c3c3c66999966,
64'h6996699666999966,
64'h0ff00ff00f0ff0f0,
64'h6699996600000000,
64'hcccccccc0ff00ff0,
64'h5555aaaac3c33c3c,
64'h3cc3c33cc33cc33c,
64'hf0f0f0f099996666,
64'h999966663cc3c33c,
64'h0f0ff0f000000000,
64'hcc3333cc0ff00ff0,
64'h66999966ff00ff00,
64'h6699996696969696,
64'hcc3333cc69966996,
64'h0000000066666666,
64'ha5a55a5a5555aaaa,
64'h3cc3c33c00000000,
64'h66666666aa5555aa,
64'h96969696aaaaaaaa,
64'h66999966aa5555aa,
64'h5aa5a55a69966996,
64'h5aa5a55a69699696,
64'h0000000099669966,
64'h99996666f00f0ff0,
64'hcc3333cc66999966,
64'hf0f0f0f0ffff0000,
64'h0000000000ffff00,
64'h699669963333cccc,
64'hc33cc33cffff0000,
64'hcc3333cc33cc33cc,
64'ha5a55a5a5aa5a55a,
64'h3333cccc00ffff00,
64'h55aa55aa55aa55aa,
64'hcc3333cccc3333cc,
64'h66666666ff00ff00,
64'h699669963c3c3c3c,
64'haa5555aa66999966,
64'hffff000066999966,
64'haaaaaaaac3c33c3c,
64'hffff0000ffff0000,
64'haa5555aac33cc33c,
64'hf00f0ff099669966,
64'h99669966ff00ff00,
64'h6996699666666666,
64'haa5555aacc3333cc,
64'hf0f0f0f03333cccc,
64'h33cc33ccf00f0ff0,
64'h0f0ff0f05555aaaa,
64'h0ff00ff0c33cc33c,
64'hcc3333cc3c3c3c3c,
64'h5aa5a55a5555aaaa,
64'h0000000069699696,
64'hcc3333cc5a5a5a5a,
64'h00ffff00f0f0f0f0,
64'h0ff00ff0aaaaaaaa,
64'hc3c33c3cc33cc33c,
64'hf0f0f0f00f0ff0f0,
64'h33cc33cc5a5a5a5a,
64'h69966996aaaaaaaa,
64'hc33cc33c96969696,
64'ha55aa55aaa5555aa,
64'h5555aaaacccccccc,
64'h00ffff00aaaaaaaa,
64'h3333cccc00ffff00,
64'h000000005aa5a55a,
64'hcc3333cc99669966,
64'hc33cc33ccccccccc,
64'h9999666600ffff00,
64'h5a5a5a5ac3c33c3c,
64'h00000000f00f0ff0,
64'h5a5a5a5a0f0ff0f0,
64'h66999966a5a55a5a,
64'ha55aa55a96969696,
64'h3333cccc3c3c3c3c,
64'h99669966ff00ff00,
64'ha55aa55a96696996,
64'h55aa55aacccccccc,
64'h3333cccc00ffff00,
64'h5555aaaa69966996,
64'h99669966a55aa55a,
64'h3333cccc5555aaaa,
64'h69699696a55aa55a,
64'h55aa55aa69966996,
64'ha5a55a5a0f0ff0f0,
64'h6996699696969696,
64'h96969696cc3333cc,
64'h5555aaaa66666666,
64'h999966660ff00ff0,
64'hccccccccff00ff00,
64'h00ffff005555aaaa,
64'h966969965a5a5a5a,
64'h0f0ff0f066666666,
64'h6699996666999966,
64'h55aa55aa66666666,
64'h33cc33cc00000000,
64'haa5555aa3c3c3c3c,
64'haa5555aaa5a55a5a,
64'hf0f0f0f069966996,
64'h96696996c33cc33c,
64'h0ff00ff096969696,
64'hffff00003cc3c33c,
64'h00ffff0033cc33cc,
64'h66666666aaaaaaaa,
64'hc33cc33cff00ff00,
64'h5aa5a55a69699696,
64'h99996666ff00ff00,
64'h00000000cccccccc,
64'h99996666f0f0f0f0,
64'haa5555aaf0f0f0f0,
64'h0f0ff0f03333cccc,
64'haaaaaaaa33cc33cc,
64'h33cc33ccaa5555aa,
64'ha55aa55a0ff00ff0,
64'hc33cc33c0ff00ff0,
64'hffff000099669966,
64'haaaaaaaaf0f0f0f0,
64'hc3c33c3c69699696,
64'hf0f0f0f0cc3333cc,
64'h9696969696696996,
64'h5555aaaac3c33c3c,
64'h9696969600ffff00,
64'h3c3c3c3c3333cccc,
64'hf00f0ff03cc3c33c,
64'h9966996666666666,
64'h3cc3c33c3c3c3c3c,
64'h55aa55aaf00f0ff0,
64'h99669966c33cc33c,
64'h5a5a5a5a66999966,
64'hc3c33c3cc33cc33c,
64'haa5555aaf0f0f0f0,
64'h33cc33ccc33cc33c,
64'hcccccccc3c3c3c3c,
64'h3333cccca55aa55a,
64'h0000000033cc33cc,
64'hc3c33c3c5a5a5a5a,
64'haa5555aaaaaaaaaa,
64'ha55aa55a69699696,
64'h5aa5a55a96969696,
64'hff00ff005aa5a55a,
64'h9999666600ffff00,
64'ha55aa55ac33cc33c,
64'hf00f0ff033cc33cc,
64'h66666666a55aa55a,
64'h0ff00ff033cc33cc,
64'h5a5a5a5a00000000,
64'h996699660ff00ff0,
64'hcccccccc66666666,
64'h66666666ff00ff00,
64'h00ffff00f00f0ff0,
64'h33cc33cccccccccc,
64'h55aa55aaf0f0f0f0,
64'ha55aa55a66999966,
64'h666666660f0ff0f0,
64'h3c3c3c3ccccccccc,
64'h0000000066999966,
64'h9696969696969696,
64'h000000005aa5a55a,
64'h0000000096696996,
64'h99669966ffff0000,
64'hffff000066666666,
64'hc33cc33c69699696,
64'h9696969699669966,
64'hc3c33c3ca55aa55a,
64'h3cc3c33c99996666,
64'ha55aa55a5aa5a55a,
64'hf0f0f0f066999966,
64'h6969969600ffff00,
64'hcc3333cc3333cccc,
64'h0ff00ff0ff00ff00,
64'h69699696aa5555aa,
64'haaaaaaaa69699696,
64'h69699696a5a55a5a,
64'hcc3333cccccccccc,
64'hf0f0f0f05aa5a55a,
64'h00ffff000f0ff0f0,
64'h00ffff000f0ff0f0,
64'ha5a55a5a66666666,
64'h0ff00ff069699696,
64'h55aa55aaaa5555aa,
64'hccccccccc33cc33c,
64'hffff000066999966,
64'hcc3333cc69699696,
64'h99996666cc3333cc,
64'h996699660ff00ff0,
64'h3cc3c33caa5555aa,
64'h96969696cccccccc,
64'h996699665555aaaa,
64'h3333cccc33cc33cc,
64'haa5555aaa55aa55a,
64'haaaaaaaac3c33c3c,
64'hf00f0ff05a5a5a5a,
64'haa5555aaffff0000,
64'h9669699696696996,
64'h696996963cc3c33c,
64'h0ff00ff0ffff0000,
64'h0000000000000000,
64'h6666666699669966,
64'hf0f0f0f05aa5a55a,
64'hc33cc33c0f0ff0f0,
64'h9696969699669966,
64'h66666666c3c33c3c,
64'h5a5a5a5affff0000,
64'h6666666600ffff00,
64'h6996699696696996,
64'h6969969633cc33cc,
64'h00ffff0066666666,
64'h00ffff005555aaaa,
64'hcc3333cc99669966,
64'haaaaaaaac3c33c3c,
64'h55aa55aa0f0ff0f0,
64'h996699665a5a5a5a,
64'hc3c33c3cc3c33c3c,
64'h5a5a5a5a33cc33cc,
64'h99996666ff00ff00,
64'haa5555aa5555aaaa,
64'h69699696cc3333cc,
64'hcccccccc5a5a5a5a,
64'hf00f0ff05a5a5a5a,
64'h966969960f0ff0f0,
64'h55aa55aac33cc33c,
64'h6969969696696996,
64'h6666666696696996,
64'h00ffff00a55aa55a,
64'ha5a55a5a00ffff00,
64'h3c3c3c3ccccccccc,
64'h3cc3c33ccc3333cc,
64'h69966996cc3333cc,
64'h0f0ff0f0cccccccc,
64'h666666665aa5a55a,
64'h69966996a55aa55a,
64'h3333cccccc3333cc,
64'h0f0ff0f05a5a5a5a,
64'ha5a55a5ac33cc33c,
64'h000000005aa5a55a,
64'hc33cc33c69966996,
64'h0f0ff0f05a5a5a5a,
64'h6996699666999966,
64'h5a5a5a5a5a5a5a5a,
64'h9669699696696996,
64'haa5555aa69966996,
64'haaaaaaaa99996666,
64'h0f0ff0f0ffff0000,
64'h00000000c3c33c3c,
64'hc33cc33c00000000,
64'haaaaaaaa00000000,
64'h999966665aa5a55a,
64'h666666660ff00ff0,
64'hc33cc33c55aa55aa,
64'h0ff00ff00f0ff0f0,
64'hcc3333ccf00f0ff0,
64'hffff0000f00f0ff0,
64'ha55aa55a00000000,
64'h55aa55aacccccccc,
64'h5aa5a55aaa5555aa,
64'h3c3c3c3c3cc3c33c,
64'h3c3c3c3c96696996,
64'h3cc3c33cffff0000,
64'ha5a55a5a33cc33cc,
64'hf0f0f0f05aa5a55a,
64'h6666666600ffff00,
64'h5aa5a55aa55aa55a,
64'h3333cccc99996666,
64'h3333cccca55aa55a,
64'h5a5a5a5aaa5555aa,
64'hc33cc33c0ff00ff0,
64'h669999663333cccc,
64'hffff00005a5a5a5a,
64'h0f0ff0f0cccccccc,
64'h96969696ffff0000,
64'h5555aaaa66999966,
64'h6996699669699696,
64'h33cc33ccf0f0f0f0,
64'hccccccccffff0000,
64'h66999966a55aa55a,
64'ha55aa55aaa5555aa,
64'h9999666655aa55aa,
64'h9669699699669966,
64'hffff000069966996,
64'h996699660ff00ff0,
64'h66999966ffff0000,
64'h33cc33cc3cc3c33c,
64'h0ff00ff05a5a5a5a,
64'haaaaaaaaffff0000,
64'h9999666696696996,
64'hff00ff00cc3333cc,
64'h3cc3c33ccccccccc,
64'ha55aa55a66999966,
64'hff00ff003cc3c33c,
64'h0f0ff0f0ff00ff00,
64'h6969969669966996,
64'haaaaaaaa0f0ff0f0,
64'hc3c33c3c96969696,
64'h0000000000ffff00,
64'h5aa5a55affff0000,
64'h00000000cccccccc,
64'h5aa5a55a99669966,
64'hcccccccc3c3c3c3c,
64'h5555aaaac3c33c3c,
64'h5a5a5a5a96969696,
64'h9999666600000000,
64'h3333cccc0ff00ff0,
64'h9669699633cc33cc,
64'h6666666696696996,
64'haaaaaaaaf00f0ff0,
64'h5a5a5a5ac33cc33c,
64'hc33cc33cf00f0ff0,
64'ha55aa55aa5a55a5a,
64'h3333cccccccccccc,
64'h3cc3c33cffff0000,
64'h33cc33ccc33cc33c,
64'h55aa55aa5555aaaa,
64'hffff0000f0f0f0f0,
64'hccccccccff00ff00,
64'h66999966ff00ff00,
64'haaaaaaaaf0f0f0f0,
64'h96969696a5a55a5a,
64'haaaaaaaa3333cccc,
64'hff00ff00aa5555aa,
64'h5a5a5a5a00ffff00,
64'h00ffff00c3c33c3c,
64'ha5a55a5aff00ff00,
64'hf0f0f0f0c33cc33c,
64'h96969696a5a55a5a,
64'h6699996696696996,
64'h5aa5a55aa55aa55a,
64'hcccccccc5555aaaa,
64'h5aa5a55a5a5a5a5a,
64'h5aa5a55a5aa5a55a,
64'h33cc33cc96969696,
64'h669999660ff00ff0,
64'h9669699600ffff00,
64'hc33cc33c5aa5a55a,
64'h69699696c3c33c3c,
64'hcc3333cc5aa5a55a,
64'hc33cc33cff00ff00,
64'h5aa5a55af00f0ff0,
64'h00ffff000ff00ff0,
64'hff00ff00cc3333cc,
64'h669999660f0ff0f0,
64'h00ffff0033cc33cc,
64'haa5555aacccccccc,
64'haa5555aac33cc33c,
64'h0f0ff0f069966996,
64'h3cc3c33ccc3333cc,
64'hf00f0ff05555aaaa,
64'h33cc33cc5aa5a55a,
64'h5a5a5a5a0f0ff0f0,
64'h99996666cc3333cc,
64'hcccccccc0f0ff0f0,
64'h3cc3c33c00000000,
64'hc3c33c3c00ffff00,
64'hf00f0ff03c3c3c3c,
64'h00000000ffff0000,
64'h0000000000ffff00,
64'ha55aa55a5a5a5a5a,
64'h69699696ff00ff00,
64'h3333ccccc3c33c3c,
64'hffff000055aa55aa,
64'h5a5a5a5a5a5a5a5a,
64'h5a5a5a5ac3c33c3c,
64'h00ffff0069966996,
64'h69966996cc3333cc,
64'hcc3333cc96696996,
64'h55aa55aaaaaaaaaa,
64'haaaaaaaa96969696,
64'hcc3333ccc33cc33c,
64'h0000000069699696,
64'h66999966cc3333cc,
64'h969696963c3c3c3c,
64'h5aa5a55a66999966,
64'h9999666669699696,
64'haa5555aa5555aaaa,
64'hf0f0f0f05a5a5a5a,
64'hf00f0ff05555aaaa,
64'h966969963333cccc,
64'h5555aaaa69966996,
64'haaaaaaaa99669966,
64'h3cc3c33c5a5a5a5a,
64'h0ff00ff0cc3333cc,
64'h33cc33cc55aa55aa,
64'h00ffff0055aa55aa,
64'hcccccccc96969696,
64'h3cc3c33cc33cc33c,
64'hf00f0ff099996666,
64'h696996965aa5a55a,
64'h5aa5a55ac3c33c3c,
64'h6666666669966996,
64'hff00ff00a5a55a5a,
64'hccccccccaa5555aa,
64'h5a5a5a5a3333cccc,
64'h5aa5a55a5a5a5a5a,
64'h99996666cccccccc,
64'h3c3c3c3ca5a55a5a,
64'h3c3c3c3ccc3333cc,
64'haa5555aa0ff00ff0,
64'h0f0ff0f099669966,
64'h00ffff0000000000,
64'h9669699696696996,
64'hffff00005aa5a55a,
64'hf0f0f0f0aaaaaaaa,
64'haaaaaaaaaaaaaaaa,
64'h96969696c3c33c3c,
64'h3cc3c33ccc3333cc,
64'h3c3c3c3c55aa55aa,
64'h9696969669699696,
64'h5555aaaa0ff00ff0,
64'h3c3c3c3caaaaaaaa,
64'h969696965555aaaa,
64'h6996699696696996,
64'h5555aaaaa5a55a5a,
64'hf0f0f0f03c3c3c3c,
64'h69699696cccccccc,
64'h6969969669699696,
64'h0f0ff0f00ff00ff0,
64'h3cc3c33c55aa55aa,
64'h9669699699669966,
64'h969696960ff00ff0,
64'h96969696a5a55a5a,
64'h99996666ffff0000,
64'h66666666cccccccc,
64'ha55aa55aa5a55a5a,
64'hffff000099669966,
64'h9999666633cc33cc,
64'ha5a55a5aff00ff00,
64'h669999665aa5a55a,
64'h999966663cc3c33c,
64'haa5555aa96696996,
64'h6996699666999966,
64'hffff0000ffff0000,
64'h5aa5a55a5a5a5a5a,
64'haa5555aa0f0ff0f0,
64'h99669966a5a55a5a,
64'h5aa5a55a5a5a5a5a,
64'hcccccccccc3333cc,
64'hf0f0f0f066999966,
64'h966969960f0ff0f0,
64'h5aa5a55a99669966,
64'h00000000f00f0ff0,
64'h5aa5a55acc3333cc,
64'h3c3c3c3c96696996,
64'h6969969633cc33cc,
64'ha5a55a5ac3c33c3c,
64'hf00f0ff099669966,
64'ha5a55a5a3cc3c33c,
64'ha55aa55a96696996,
64'hf00f0ff03c3c3c3c,
64'hc33cc33caaaaaaaa,
64'h00000000a55aa55a,
64'h5555aaaaaaaaaaaa,
64'h6666666600000000,
64'h3c3c3c3ccc3333cc,
64'h5aa5a55aaa5555aa,
64'h5a5a5a5a3333cccc,
64'h33cc33ccff00ff00,
64'hf00f0ff0aa5555aa,
64'h00ffff00aa5555aa,
64'hccccccccaaaaaaaa,
64'h99996666f0f0f0f0,
64'h3cc3c33c3333cccc,
64'h966969965aa5a55a,
64'h5555aaaa96696996,
64'h66666666aaaaaaaa,
64'h33cc33cca5a55a5a,
64'hf00f0ff0cc3333cc,
64'hf00f0ff05555aaaa,
64'h9966996666999966,
64'h3cc3c33c3c3c3c3c,
64'h6666666666999966,
64'hffff00003333cccc,
64'hc33cc33c55aa55aa,
64'h69699696f0f0f0f0,
64'h9999666699669966,
64'h0ff00ff0f0f0f0f0,
64'ha55aa55a00000000,
64'h3333cccc69699696,
64'hf0f0f0f069966996,
64'h6666666655aa55aa,
64'h0000000000000000,
64'h3c3c3c3c66999966,
64'hc3c33c3c3333cccc,
64'h9669699699996666,
64'hc3c33c3cc3c33c3c,
64'h33cc33cc3cc3c33c,
64'h00ffff0000ffff00,
64'hcc3333cc00000000,
64'h5a5a5a5a5aa5a55a,
64'h3c3c3c3c99669966,
64'h9696969600000000,
64'hc3c33c3c96696996,
64'hc33cc33ca5a55a5a,
64'h3c3c3c3c5a5a5a5a,
64'haa5555aac3c33c3c,
64'h996699665aa5a55a,
64'hc3c33c3c5555aaaa,
64'h969696963cc3c33c,
64'h0ff00ff0ff00ff00,
64'h00ffff0069966996,
64'h3c3c3c3cffff0000,
64'hccccccccaaaaaaaa,
64'h5555aaaa5a5a5a5a,
64'h00ffff00c3c33c3c,
64'hc33cc33c0ff00ff0,
64'hf0f0f0f00ff00ff0,
64'h5aa5a55a69966996,
64'haaaaaaaa00000000,
64'h5a5a5a5a00ffff00,
64'h999966660f0ff0f0,
64'ha55aa55a3cc3c33c,
64'h5aa5a55aaa5555aa,
64'hc3c33c3c5aa5a55a,
64'h3333cccc00ffff00,
64'h3c3c3c3c99669966,
64'h5555aaaa5a5a5a5a,
64'h9669699600000000,
64'h5a5a5a5a5aa5a55a,
64'hf00f0ff0cccccccc,
64'h5555aaaa55aa55aa,
64'haaaaaaaaffff0000,
64'h3cc3c33cffff0000,
64'h99669966ff00ff00,
64'h33cc33cc33cc33cc,
64'h696996965a5a5a5a,
64'hcccccccc99996666,
64'h999966665555aaaa,
64'hff00ff00a55aa55a,
64'h5aa5a55a5555aaaa,
64'haaaaaaaaf00f0ff0,
64'h0000000033cc33cc,
64'h6666666696696996,
64'hf0f0f0f066999966,
64'hff00ff00cccccccc,
64'h9966996699669966,
64'h3cc3c33ccc3333cc,
64'hff00ff0069966996,
64'h5555aaaa00ffff00,
64'h99996666ffff0000,
64'h5a5a5a5a66999966,
64'h99996666a55aa55a,
64'h6666666666999966,
64'h000000005555aaaa,
64'h3333cccc00ffff00,
64'ha55aa55aaa5555aa,
64'h5aa5a55a0f0ff0f0,
64'h0ff00ff055aa55aa,
64'h5a5a5a5aa5a55a5a,
64'haa5555aaf0f0f0f0,
64'h5555aaaaf00f0ff0,
64'h969696963cc3c33c,
64'h3333cccc0f0ff0f0,
64'h6666666666666666,
64'hf0f0f0f066999966,
64'h6969969655aa55aa,
64'h3333cccca5a55a5a,
64'h9669699655aa55aa,
64'hff00ff00aaaaaaaa,
64'ha55aa55affff0000,
64'haaaaaaaaa55aa55a,
64'h9696969600000000,
64'hffff00005555aaaa,
64'hcccccccc99669966,
64'h99669966ffff0000,
64'ha55aa55a0ff00ff0,
64'h6969969699996666,
64'hcccccccc33cc33cc,
64'h699669960ff00ff0,
64'h3c3c3c3c96696996,
64'hffff00000f0ff0f0,
64'hc33cc33c96696996,
64'h0ff00ff066666666,
64'h66666666c33cc33c,
64'h99996666f00f0ff0,
64'h69966996c33cc33c,
64'haaaaaaaaa5a55a5a,
64'ha5a55a5aa55aa55a,
64'hf00f0ff0c3c33c3c,
64'hf00f0ff069966996,
64'hf0f0f0f066666666,
64'h00ffff0099669966,
64'h5aa5a55acccccccc,
64'hc33cc33c5a5a5a5a,
64'h5555aaaa96696996,
64'h0ff00ff0c3c33c3c,
64'h6969969633cc33cc,
64'hf00f0ff00f0ff0f0,
64'hc33cc33c99996666,
64'haa5555aa3333cccc,
64'h0ff00ff0c33cc33c,
64'h66999966f00f0ff0,
64'h696996963c3c3c3c,
64'hf00f0ff066999966,
64'h3c3c3c3ca55aa55a,
64'h5555aaaa96696996,
64'h9669699633cc33cc,
64'h5555aaaa99996666,
64'h999966665a5a5a5a,
64'hff00ff0099669966,
64'hccccccccf0f0f0f0,
64'h6996699633cc33cc,
64'haa5555aaa5a55a5a,
64'hff00ff00aa5555aa,
64'h5a5a5a5ac3c33c3c,
64'hcc3333cc00000000,
64'h966969963cc3c33c,
64'h3cc3c33c66999966,
64'h0f0ff0f066666666,
64'h66666666cccccccc,
64'h699669960ff00ff0,
64'h33cc33cca5a55a5a,
64'h6969969699996666,
64'h96969696c33cc33c,
64'ha5a55a5aaa5555aa,
64'haaaaaaaacccccccc,
64'h69966996cccccccc,
64'h6996699696696996,
64'h5aa5a55a99669966,
64'hf00f0ff0a55aa55a,
64'hff00ff00f0f0f0f0,
64'ha55aa55ac33cc33c,
64'h3cc3c33caa5555aa,
64'h5555aaaa3333cccc,
64'hc3c33c3cc3c33c3c,
64'hf0f0f0f000ffff00,
64'hcccccccc33cc33cc,
64'h99996666aaaaaaaa,
64'h696996965a5a5a5a,
64'h00ffff0033cc33cc,
64'ha5a55a5a69699696,
64'h0ff00ff00f0ff0f0,
64'haaaaaaaaffff0000,
64'h96696996cc3333cc,
64'hcc3333cc5aa5a55a,
64'ha55aa55a96696996,
64'h0000000069699696,
64'h66999966aaaaaaaa,
64'h9966996699669966,
64'hc3c33c3cff00ff00,
64'h6666666699669966,
64'h6996699699669966,
64'h000000000f0ff0f0,
64'h3333cccc69699696,
64'h5a5a5a5a55aa55aa,
64'h6996699669699696,
64'h33cc33cc00ffff00,
64'h3c3c3c3ca5a55a5a,
64'h6969969696696996,
64'h5555aaaaa5a55a5a,
64'haaaaaaaa0ff00ff0,
64'h6996699669699696,
64'h00000000f00f0ff0,
64'h5a5a5a5a96696996,
64'h96969696a55aa55a,
64'h66999966cccccccc,
64'haaaaaaaacc3333cc,
64'h69966996cccccccc,
64'h3c3c3c3c00000000,
64'h0ff00ff00f0ff0f0,
64'h0000000099996666,
64'h3333cccc5a5a5a5a,
64'h3c3c3c3c5555aaaa,
64'hffff00003333cccc,
64'hff00ff0099996666,
64'hf00f0ff066666666,
64'h96969696ff00ff00,
64'haa5555aaf0f0f0f0,
64'ha55aa55a66999966,
64'h3cc3c33c96696996,
64'h00ffff0066666666,
64'ha5a55a5a33cc33cc,
64'ha55aa55aa5a55a5a,
64'h6666666666666666,
64'h3c3c3c3c69699696,
64'h96969696a55aa55a,
64'haaaaaaaac3c33c3c,
64'h669999665a5a5a5a,
64'h6996699666666666,
64'hc33cc33cff00ff00,
64'h96969696c3c33c3c,
64'haa5555aaff00ff00,
64'hcc3333cc00000000,
64'hf0f0f0f0c33cc33c,
64'h55aa55aa96696996,
64'h3c3c3c3c3333cccc,
64'h0000000000000000,
64'h0ff00ff0c3c33c3c,
64'h0ff00ff05a5a5a5a,
64'h9669699696969696,
64'ha55aa55aa55aa55a,
64'ha5a55a5a5aa5a55a,
64'hffff00005555aaaa,
64'ha5a55a5aaaaaaaaa,
64'h99669966cc3333cc,
64'h0ff00ff069699696,
64'hc33cc33c00000000,
64'h0ff00ff03cc3c33c,
64'h5aa5a55a99669966,
64'h0ff00ff099669966,
64'h3333cccc0ff00ff0,
64'h6969969666999966,
64'h0ff00ff066666666,
64'h699669965aa5a55a,
64'h00ffff005555aaaa,
64'hffff00003cc3c33c,
64'ha55aa55a00000000,
64'hf0f0f0f066666666,
64'hcccccccc33cc33cc,
64'h5555aaaa0ff00ff0,
64'h5aa5a55aaa5555aa,
64'hff00ff0000ffff00,
64'hcc3333cc3cc3c33c,
64'h6666666600000000,
64'h33cc33ccffff0000,
64'h3c3c3c3c55aa55aa,
64'h669999665aa5a55a,
64'hcc3333cc99996666,
64'ha55aa55a66999966,
64'h5a5a5a5a5555aaaa,
64'ha55aa55a69699696,
64'hcccccccc33cc33cc,
64'h9669699600000000,
64'h99669966cc3333cc,
64'h00ffff005a5a5a5a,
64'h666666663333cccc,
64'h6666666600000000,
64'hf00f0ff0aaaaaaaa,
64'h696996965555aaaa,
64'h0f0ff0f00f0ff0f0,
64'hc33cc33c33cc33cc,
64'h5a5a5a5a3c3c3c3c,
64'h3c3c3c3c66666666,
64'h5555aaaa66999966,
64'hcc3333cccccccccc,
64'h66666666aa5555aa,
64'h00000000a5a55a5a,
64'h3c3c3c3c3cc3c33c,
64'hff00ff0069699696,
64'hffff00005a5a5a5a,
64'hc3c33c3cc3c33c3c,
64'hf00f0ff00f0ff0f0,
64'h5555aaaa96696996,
64'hccccccccffff0000,
64'h96969696aaaaaaaa,
64'h9966996669699696,
64'h3c3c3c3c66999966,
64'h96969696c3c33c3c,
64'h0000000066666666,
64'hf0f0f0f05555aaaa,
64'h6699996699996666,
64'hcc3333cc55aa55aa,
64'haa5555aa99996666,
64'h33cc33cc33cc33cc,
64'h3333cccc55aa55aa,
64'h6666666600ffff00,
64'h699669965aa5a55a,
64'hf0f0f0f055aa55aa,
64'h9696969696969696,
64'hff00ff00c3c33c3c,
64'hc33cc33c99996666,
64'h5a5a5a5a33cc33cc,
64'h9669699699996666,
64'h5555aaaacccccccc,
64'hcc3333cc00000000,
64'hcccccccc66999966,
64'hc33cc33c00000000,
64'h00000000cccccccc,
64'h5a5a5a5a69699696,
64'hc3c33c3c00000000,
64'hcc3333ccaa5555aa,
64'hc33cc33c3c3c3c3c,
64'h5a5a5a5aa5a55a5a,
64'h3cc3c33c00ffff00,
64'h0ff00ff03cc3c33c,
64'h0000000055aa55aa,
64'h5aa5a55a96696996,
64'h00ffff0096969696,
64'h3c3c3c3cf00f0ff0,
64'h3c3c3c3c00ffff00,
64'h966969965aa5a55a,
64'hcccccccc33cc33cc,
64'h33cc33cc66999966,
64'haa5555aa0ff00ff0,
64'haa5555aa96696996,
64'h55aa55aa3c3c3c3c,
64'hffff0000c3c33c3c,
64'h66999966f0f0f0f0,
64'h5aa5a55a33cc33cc,
64'hcccccccc3cc3c33c,
64'haa5555aaa55aa55a,
64'hc33cc33ca5a55a5a,
64'haa5555aaff00ff00,
64'h5aa5a55a96969696,
64'h3333cccc5a5a5a5a,
64'haa5555aa5aa5a55a,
64'hc3c33c3c00ffff00,
64'h69966996a55aa55a,
64'haa5555aac3c33c3c,
64'ha55aa55a66999966,
64'hcccccccc3cc3c33c,
64'h96696996a5a55a5a,
64'h666666663c3c3c3c,
64'h9696969699669966,
64'h5555aaaac3c33c3c,
64'hf0f0f0f0ff00ff00,
64'h3cc3c33c0f0ff0f0,
64'h3333cccc33cc33cc,
64'h5555aaaa99996666,
64'h33cc33cca55aa55a,
64'h0f0ff0f0aaaaaaaa,
64'h96696996f00f0ff0,
64'h5aa5a55a69699696,
64'h55aa55aa96969696,
64'h96969696f0f0f0f0,
64'h3cc3c33c00ffff00,
64'h0f0ff0f033cc33cc,
64'hc33cc33c96969696,
64'h699669965aa5a55a,
64'h33cc33cc3333cccc,
64'h666666665a5a5a5a,
64'h3cc3c33cf0f0f0f0,
64'h3cc3c33c3cc3c33c,
64'hcc3333cc69699696,
64'haa5555aacc3333cc,
64'h5555aaaaff00ff00,
64'hcc3333ccf00f0ff0,
64'hf00f0ff03333cccc,
64'h666666665a5a5a5a,
64'ha55aa55aa55aa55a,
64'h55aa55aa5555aaaa,
64'hf0f0f0f0a5a55a5a,
64'h3c3c3c3ccccccccc,
64'h6996699633cc33cc,
64'h5555aaaa0f0ff0f0,
64'h99669966c33cc33c,
64'haa5555aa55aa55aa,
64'hccccccccaaaaaaaa,
64'h3cc3c33ca5a55a5a,
64'ha5a55a5a66999966,
64'h6699996696696996,
64'h0000000069966996,
64'hc3c33c3c66666666,
64'h69699696c3c33c3c,
64'h0ff00ff0ffff0000,
64'h96969696c3c33c3c,
64'h3cc3c33cc3c33c3c,
64'h00000000ff00ff00,
64'hf0f0f0f069966996,
64'h9966996699996666,
64'h3cc3c33cc33cc33c,
64'h0f0ff0f05555aaaa,
64'h0ff00ff099669966,
64'hc33cc33c96696996,
64'h6666666699669966,
64'h66666666aa5555aa,
64'h3cc3c33cc33cc33c,
64'h00000000aa5555aa,
64'h33cc33cc96696996,
64'hc33cc33c66999966,
64'hc3c33c3cf0f0f0f0,
64'h666666660f0ff0f0,
64'h3cc3c33c5a5a5a5a,
64'h0ff00ff000000000,
64'h00ffff00ff00ff00,
64'h0000000096969696,
64'hf0f0f0f099669966,
64'ha55aa55acccccccc,
64'h000000005a5a5a5a,
64'h5555aaaa96969696,
64'h00ffff0096969696,
64'h69966996ffff0000,
64'h3333ccccff00ff00,
64'h66999966c3c33c3c,
64'hf00f0ff096696996,
64'h5555aaaa96969696,
64'h996699660f0ff0f0,
64'h6699996633cc33cc,
64'h3c3c3c3c96969696,
64'h0ff00ff0c33cc33c,
64'hc33cc33c66999966,
64'hcccccccc0ff00ff0,
64'hc3c33c3c99669966,
64'h699669963c3c3c3c,
64'hf00f0ff0ffff0000,
64'hc33cc33c0ff00ff0,
64'h3333cccc5555aaaa,
64'ha5a55a5a00000000,
64'h55aa55aaf00f0ff0,
64'h3333cccc3cc3c33c,
64'h0ff00ff05a5a5a5a,
64'h00000000aaaaaaaa,
64'h00ffff000ff00ff0,
64'h00ffff0099669966,
64'h3cc3c33cc33cc33c,
64'h66999966cc3333cc,
64'h33cc33cccc3333cc,
64'haaaaaaaa66666666,
64'h9966996666666666,
64'h696996960f0ff0f0,
64'h00ffff0069966996,
64'hf00f0ff0aaaaaaaa,
64'h00ffff00f00f0ff0,
64'hcc3333cc69699696,
64'haa5555aac3c33c3c,
64'hf0f0f0f000ffff00,
64'h69966996c3c33c3c,
64'haa5555aa96969696,
64'h3cc3c33ccc3333cc,
64'hffff000066666666,
64'haaaaaaaa5aa5a55a,
64'h66999966aaaaaaaa,
64'hff00ff003c3c3c3c,
64'hf0f0f0f00f0ff0f0,
64'hcccccccc00ffff00,
64'h669999663333cccc,
64'h5555aaaa5555aaaa,
64'h0f0ff0f05aa5a55a,
64'h96969696aaaaaaaa,
64'h0f0ff0f000000000,
64'h0ff00ff099996666,
64'hc3c33c3ccc3333cc,
64'ha5a55a5a96969696,
64'h6699996669699696,
64'h33cc33cc66666666,
64'hcc3333cc69966996,
64'hf0f0f0f0a5a55a5a,
64'h3cc3c33c00000000,
64'h696996960f0ff0f0,
64'hffff000099669966,
64'h96969696f0f0f0f0,
64'h3c3c3c3caaaaaaaa,
64'h00ffff00cccccccc,
64'h69966996cccccccc,
64'h55aa55aa55aa55aa,
64'h5aa5a55aa5a55a5a,
64'h33cc33cc0ff00ff0,
64'h0ff00ff03c3c3c3c,
64'hccccccccc3c33c3c,
64'ha5a55a5a5a5a5a5a,
64'h969696963333cccc,
64'h0000000099669966,
64'h0ff00ff05aa5a55a,
64'hffff000069966996,
64'h0000000099669966,
64'ha55aa55a0ff00ff0,
64'haa5555aa55aa55aa,
64'h6666666696696996,
64'h5a5a5a5aaaaaaaaa,
64'hc33cc33c66666666,
64'hc3c33c3cc33cc33c,
64'h0ff00ff069699696,
64'hc33cc33ca55aa55a,
64'h0000000096969696,
64'hff00ff00cccccccc,
64'hc3c33c3c96969696,
64'ha5a55a5a99996666,
64'h999966663c3c3c3c,
64'ha5a55a5aa5a55a5a,
64'hf0f0f0f03333cccc,
64'h96969696ffff0000,
64'h3cc3c33c66999966,
64'hff00ff0099996666,
64'hc33cc33cc33cc33c,
64'hffff00000ff00ff0,
64'hf00f0ff096969696,
64'h33cc33cca5a55a5a,
64'h3cc3c33c3c3c3c3c,
64'h666666665a5a5a5a,
64'ha5a55a5a00000000,
64'h5a5a5a5ac3c33c3c,
64'hf00f0ff0aaaaaaaa,
64'h00000000f0f0f0f0,
64'h33cc33ccc33cc33c,
64'h0ff00ff0aaaaaaaa,
64'ha5a55a5a3333cccc,
64'h5aa5a55aa55aa55a,
64'h33cc33cc33cc33cc,
64'hf00f0ff05555aaaa,
64'haa5555aa5aa5a55a,
64'h0000000099996666,
64'hcc3333cc3cc3c33c,
64'h5555aaaa69966996,
64'ha55aa55a00ffff00,
64'h0ff00ff05555aaaa,
64'h3cc3c33c66999966,
64'h5a5a5a5aa5a55a5a,
64'h0f0ff0f0c3c33c3c,
64'h3333ccccaa5555aa,
64'h999966663cc3c33c,
64'h99996666a55aa55a,
64'h000000000ff00ff0,
64'h6969969655aa55aa,
64'h669999660f0ff0f0,
64'h5a5a5a5af00f0ff0,
64'h3333cccc66999966,
64'h5aa5a55a33cc33cc,
64'h3333cccc5555aaaa,
64'h66999966c33cc33c,
64'h5a5a5a5a33cc33cc,
64'h99996666cc3333cc,
64'ha55aa55a5555aaaa,
64'h9669699666999966,
64'h3333cccc0ff00ff0,
64'h6699996669699696,
64'hf0f0f0f05aa5a55a,
64'h3cc3c33c99669966,
64'h96969696a55aa55a,
64'hc33cc33cc3c33c3c,
64'hcccccccc0ff00ff0,
64'h55aa55aa5555aaaa,
64'hf00f0ff0ff00ff00,
64'h5a5a5a5aa5a55a5a,
64'h666666663c3c3c3c,
64'ha5a55a5a66999966,
64'hff00ff00cccccccc,
64'h9669699600ffff00,
64'h6699996669966996,
64'h9999666669966996,
64'hc33cc33cff00ff00,
64'hf00f0ff0ffff0000,
64'h55aa55aaa5a55a5a,
64'h5aa5a55ac33cc33c,
64'h3cc3c33ccc3333cc,
64'h0f0ff0f05a5a5a5a,
64'h3c3c3c3c99669966,
64'hf00f0ff0ff00ff00,
64'h5aa5a55af00f0ff0,
64'ha5a55a5a69966996,
64'h99996666a5a55a5a,
64'h666666665555aaaa,
64'ha5a55a5a00ffff00,
64'haa5555aa5a5a5a5a,
64'h9696969699669966,
64'hcc3333cccc3333cc,
64'h3333cccccccccccc,
64'hff00ff0099669966,
64'h0ff00ff05a5a5a5a,
64'h3cc3c33c0f0ff0f0,
64'hccccccccff00ff00,
64'h696996965aa5a55a,
64'h3333cccc3333cccc,
64'h5a5a5a5acccccccc,
64'hf00f0ff033cc33cc,
64'h9966996669699696,
64'h6969969696696996,
64'haaaaaaaa96696996,
64'h0ff00ff03c3c3c3c,
64'h699669960ff00ff0,
64'haa5555aaaaaaaaaa,
64'hc33cc33ca55aa55a,
64'hf00f0ff0a55aa55a,
64'haaaaaaaa5555aaaa,
64'hff00ff003cc3c33c,
64'hc3c33c3c3c3c3c3c,
64'hf00f0ff05aa5a55a,
64'h55aa55aacccccccc,
64'haa5555aa69699696,
64'hf00f0ff03cc3c33c,
64'h3c3c3c3c69699696,
64'h3c3c3c3c3333cccc,
64'hf00f0ff05aa5a55a,
64'haaaaaaaa3333cccc,
64'h0f0ff0f096696996,
64'hf00f0ff069699696,
64'h0ff00ff055aa55aa,
64'h96969696ff00ff00,
64'hf00f0ff099669966,
64'haa5555aa00000000,
64'hffff0000ffff0000,
64'haaaaaaaac33cc33c,
64'hff00ff00c3c33c3c,
64'hcc3333ccf0f0f0f0,
64'h0000000033cc33cc,
64'hccccccccc33cc33c,
64'h5555aaaac33cc33c,
64'h9669699600000000,
64'hf0f0f0f05555aaaa,
64'h696996960ff00ff0,
64'haa5555aa96696996,
64'h6666666669966996,
64'h69699696ff00ff00,
64'hc3c33c3ca5a55a5a,
64'ha55aa55ac33cc33c,
64'h00ffff00f00f0ff0,
64'hf00f0ff0c3c33c3c,
64'hf0f0f0f0aa5555aa,
64'h0ff00ff0c3c33c3c,
64'h699669960ff00ff0,
64'h00ffff0000000000,
64'h5aa5a55aaa5555aa,
64'hf0f0f0f0cccccccc,
64'h99669966aaaaaaaa,
64'h9999666600ffff00,
64'hf0f0f0f05aa5a55a,
64'haa5555aa99669966,
64'h00000000cccccccc,
64'hffff000000ffff00,
64'h5555aaaac3c33c3c,
64'h5aa5a55af00f0ff0,
64'h696996960f0ff0f0,
64'ha5a55a5aa5a55a5a,
64'hcccccccc96969696,
64'hc3c33c3c3c3c3c3c,
64'hc33cc33cff00ff00,
64'h5555aaaa96696996,
64'haa5555aacccccccc,
64'h5555aaaa00ffff00,
64'ha5a55a5a69966996,
64'h99996666a55aa55a,
64'h55aa55aa5555aaaa,
64'h3cc3c33ca55aa55a,
64'h3333cccc69966996,
64'h5aa5a55a0f0ff0f0,
64'haaaaaaaa96969696,
64'h66666666cc3333cc,
64'hc3c33c3c66666666,
64'h5555aaaa0ff00ff0,
64'hff00ff00ff00ff00,
64'hf0f0f0f05555aaaa,
64'hc3c33c3c5a5a5a5a,
64'h6666666666666666,
64'h55aa55aa66999966,
64'h6996699666666666,
64'hff00ff0000000000,
64'haa5555aa3c3c3c3c,
64'h0ff00ff0a5a55a5a,
64'h9966996669966996,
64'h69699696c33cc33c,
64'ha5a55a5a96969696,
64'h0f0ff0f03cc3c33c,
64'h55aa55aa33cc33cc,
64'hf00f0ff0aaaaaaaa,
64'h69966996ff00ff00,
64'haaaaaaaa69699696,
64'h69966996ff00ff00,
64'h0ff00ff0cccccccc,
64'hffff0000f0f0f0f0,
64'h96696996f0f0f0f0,
64'h3333cccc3333cccc,
64'hcc3333cc33cc33cc,
64'ha5a55a5aaa5555aa,
64'h00ffff000ff00ff0,
64'hf0f0f0f00ff00ff0,
64'h33cc33cc99669966,
64'h69966996f0f0f0f0,
64'h0000000069699696,
64'h00ffff00cc3333cc,
64'h0000000096696996,
64'haaaaaaaac3c33c3c,
64'hcc3333cc00ffff00,
64'h3333cccc3333cccc,
64'h969696963cc3c33c,
64'h33cc33cc66666666,
64'hf00f0ff03c3c3c3c,
64'h0ff00ff0f00f0ff0,
64'haa5555aac33cc33c,
64'hf00f0ff066999966,
64'h00000000c33cc33c,
64'hffff0000f0f0f0f0,
64'h0ff00ff0c33cc33c,
64'h996699663c3c3c3c,
64'h96969696a55aa55a,
64'h9966996633cc33cc,
64'h55aa55aa5a5a5a5a,
64'hc33cc33caaaaaaaa,
64'hf00f0ff069699696,
64'h5555aaaa96969696,
64'hf00f0ff05aa5a55a,
64'h0000000000ffff00,
64'haa5555aac33cc33c,
64'ha5a55a5a33cc33cc,
64'hf00f0ff0a55aa55a,
64'h9696969633cc33cc,
64'h33cc33cc00000000,
64'h996699660ff00ff0,
64'h00ffff0066666666,
64'haaaaaaaaff00ff00,
64'h0f0ff0f0f00f0ff0,
64'h00ffff00cccccccc,
64'h33cc33ccf0f0f0f0,
64'h6699996666999966,
64'ha5a55a5a0f0ff0f0,
64'h00ffff00cccccccc,
64'h9999666666999966,
64'haaaaaaaa96969696,
64'h0f0ff0f05aa5a55a,
64'h6666666696696996,
64'h66999966ffff0000,
64'h00ffff0066666666,
64'hf00f0ff069699696,
64'h9966996699669966,
64'hff00ff00a55aa55a,
64'h5a5a5a5a99996666,
64'h969696965aa5a55a,
64'h9696969666999966,
64'haaaaaaaa00ffff00,
64'hc33cc33c3333cccc,
64'h69699696ff00ff00,
64'h99669966aa5555aa,
64'hf0f0f0f069699696,
64'h66999966a5a55a5a,
64'h5a5a5a5acccccccc,
64'h696996965aa5a55a,
64'h996699660f0ff0f0,
64'h3c3c3c3c0f0ff0f0,
64'h6699996666666666,
64'h3cc3c33c69699696,
64'h5a5a5a5aaa5555aa,
64'h69699696c33cc33c,
64'h55aa55aa66999966,
64'hf00f0ff069699696,
64'h69966996cc3333cc,
64'hf00f0ff00ff00ff0,
64'hf0f0f0f0aa5555aa,
64'h3333cccccccccccc,
64'h00ffff005555aaaa,
64'h9966996633cc33cc,
64'h3c3c3c3ca55aa55a,
64'h33cc33ccc3c33c3c,
64'h5555aaaa5a5a5a5a,
64'h3cc3c33cffff0000,
64'h6969969696696996,
64'h969696963cc3c33c,
64'h5aa5a55affff0000,
64'h00ffff0000000000,
64'h9999666699669966,
64'hcc3333cc5aa5a55a,
64'h5aa5a55a0f0ff0f0,
64'h55aa55aa99669966,
64'ha55aa55ac3c33c3c,
64'h00ffff00ffff0000,
64'h6699996600ffff00,
64'h9966996696696996,
64'h9696969633cc33cc,
64'h9696969666666666,
64'h33cc33cc5555aaaa,
64'h9999666699669966,
64'h69966996c3c33c3c,
64'h0f0ff0f00f0ff0f0,
64'h5a5a5a5a5a5a5a5a,
64'h5555aaaac3c33c3c,
64'h00ffff0033cc33cc,
64'hf00f0ff0ff00ff00,
64'h5a5a5a5a5555aaaa,
64'hc33cc33ccc3333cc,
64'h5a5a5a5a5a5a5a5a,
64'h996699665a5a5a5a,
64'h00ffff000f0ff0f0,
64'h69699696c33cc33c,
64'hc33cc33c96696996,
64'h6666666696696996,
64'h00ffff00a55aa55a,
64'h3cc3c33c00ffff00,
64'h3333cccccccccccc,
64'h5aa5a55acc3333cc,
64'h00ffff00cc3333cc,
64'h66666666cccccccc,
64'hffff00005aa5a55a,
64'h0ff00ff0a55aa55a,
64'haa5555aacc3333cc,
64'h999966665a5a5a5a,
64'h3333ccccc33cc33c,
64'haa5555aa5aa5a55a,
64'ha55aa55a69966996,
64'h0ff00ff05a5a5a5a,
64'h00ffff0066999966,
64'h666666665a5a5a5a,
64'hff00ff0096696996,
64'haa5555aa69966996,
64'haa5555aa99996666,
64'hc33cc33cffff0000,
64'h00ffff00c3c33c3c,
64'h9999666600000000,
64'haaaaaaaa00000000,
64'h666666665aa5a55a,
64'hffff00000ff00ff0,
64'h0f0ff0f055aa55aa,
64'haaaaaaaa0f0ff0f0,
64'hf0f0f0f0f00f0ff0,
64'hccccccccf00f0ff0,
64'h9669699600000000,
64'h55aa55aacccccccc,
64'hc33cc33caa5555aa,
64'h999966663cc3c33c,
64'h9696969696696996,
64'hc33cc33cffff0000,
64'ha55aa55a33cc33cc,
64'h669999665aa5a55a,
64'hffff000000ffff00,
64'haa5555aaa55aa55a,
64'h55aa55aa99996666,
64'h00ffff00a55aa55a,
64'hc33cc33c55aa55aa

 } ; 


wire [LUT_NUM_ONE_EQUATION*2*16-1:0]  dout_pre ;


genvar i,j;
generate
    for (i=0; i<16; i=i+1) begin : first_layer_1
    	for (j=0; j<LUT_NUM_ONE_EQUATION; j=j+1) begin : first_layer_2
    	 //   	LUT6 #(
		   	//    .INIT(POLY[i*LUT_NUM_ONE_EQUATION*64+j*64 +: 64])  // Specify LUT Contents
		   	// ) LUT6_inst (
		   	//    .O(dout_pre[i*LUT_NUM_ONE_EQUATION+j]),   // LUT general output
		   	//    .I0(din[j*6]  ), // LUT input
		   	//    .I1(din[j*6+1]), // LUT input
		   	//    .I2(din[j*6+2]), // LUT input
		   	//    .I3(din[j*6+3]), // LUT input
		   	//    .I4(din[j*6+4]), // LUT input
		   	//    .I5(din[j*6+5])  // LUT input
		   	// );
   			LUT6_2 #(
   			   .INIT(POLY[i*LUT_NUM_ONE_EQUATION*64+j*64 +: 64]) // Specify LUT Contents
   			) LUT6_2_inst (
   			   .O6(dout_pre[i*LUT_NUM_ONE_EQUATION+j]), // 1-bit LUT6 output
   			   .O5(dout_pre[i*LUT_NUM_ONE_EQUATION+j+16*LUT_NUM_ONE_EQUATION]), // 1-bit lower LUT5 output
   			   .I0(din[j*5]  ), // 1-bit LUT input
   			   .I1(din[j*5+1]), // 1-bit LUT input
   			   .I2(din[j*5+2]), // 1-bit LUT input
   			   .I3(din[j*5+3]), // 1-bit LUT input
   			   .I4(din[j*5+4]), // 1-bit LUT input
   			   .I5(1'b1)  // 1-bit LUT input (fast MUX select only available to O6 output)
   			);
    	end
    end
endgenerate






integer m,n ;
always @(posedge clk or posedge rst) begin
	if (rst == 1'b1) begin
		dout <= 'b0 ;
	end
    else begin
    	for (m=0; m<32; m=m+1) begin 
    		for (n=0; n<LUT_OUT_NUM_ONE_EQUATION; n=n+1) begin 
    			if ( n<LUT_NUM_ONE_EQUATION ) begin
    				dout[m*LUT_OUT_NUM_ONE_EQUATION+n] <= dout_pre[m*LUT_NUM_ONE_EQUATION+n];
    			end
    			else begin
    				dout[m*LUT_OUT_NUM_ONE_EQUATION+n] <= 1'b0 ;
    			end
    		end
    	end
    end
end




endmodule 

// always @(posedge clk or posedge rst) begin
// 	if (rst == 1'b1) begin
// 		dout <= 'b0 ;
// 	end
//     else begin
//        dout <= dout_pre ; 
//     end
// end