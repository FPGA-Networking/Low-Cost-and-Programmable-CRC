


module layer_1_new 
    # ( parameter  LUT_NUM_ONE_EQUATION    		  = 0 , // 171      // and thre are 32 equation
    			         LUT_OUT_NUM_ONE_EQUATION     = 0 , // 174
                   LUT_POLY                     = 0 ,                   
    	             BUS_WIDTH  		              = LUT_NUM_ONE_EQUATION*5  
        )
( 
            input	            		clk      ,   
            input	            		rst      ,   
            input      [BUS_WIDTH-1:0]    	din      ,
            output reg [LUT_OUT_NUM_ONE_EQUATION*32-1:0]       dout 				      

 ) ;






parameter  [0:LUT_NUM_ONE_EQUATION*64*16-1] POLY  = LUT_POLY ;


wire [LUT_NUM_ONE_EQUATION*2*16-1:0]  dout_pre ;


genvar i,j;
generate
    for (i=0; i<16; i=i+1) begin : first_layer_1
    	for (j=0; j<LUT_NUM_ONE_EQUATION; j=j+1) begin : first_layer_2
    	 //   	LUT6 #(
		   	//    .INIT(POLY[i*LUT_NUM_ONE_EQUATION*64+j*64 +: 64])  // Specify LUT Contents
		   	// ) LUT6_inst (
		   	//    .O(dout_pre[i*LUT_NUM_ONE_EQUATION+j]),   // LUT general output
		   	//    .I0(din[j*6]  ), // LUT input
		   	//    .I1(din[j*6+1]), // LUT input
		   	//    .I2(din[j*6+2]), // LUT input
		   	//    .I3(din[j*6+3]), // LUT input
		   	//    .I4(din[j*6+4]), // LUT input
		   	//    .I5(din[j*6+5])  // LUT input
		   	// );
(* DONT_TOUCH= "TRUE" *)  			LUT6_2 #(
   			   .INIT(POLY[i*LUT_NUM_ONE_EQUATION*64+j*64 +: 64]) // Specify LUT Contents
   			) LUT6_2_inst (
   			   .O6(dout_pre[i*LUT_NUM_ONE_EQUATION+j]), // 1-bit LUT6 output
   			   .O5(dout_pre[i*LUT_NUM_ONE_EQUATION+j+16*LUT_NUM_ONE_EQUATION]), // 1-bit lower LUT5 output
   			   .I0(din[j*5]  ), // 1-bit LUT input
   			   .I1(din[j*5+1]), // 1-bit LUT input
   			   .I2(din[j*5+2]), // 1-bit LUT input
   			   .I3(din[j*5+3]), // 1-bit LUT input
   			   .I4(din[j*5+4]), // 1-bit LUT input
   			   .I5(1'b1)  // 1-bit LUT input (fast MUX select only available to O6 output)
   			);
    	end
    end
endgenerate






// integer m,n ;
// always @(posedge clk or posedge rst) begin
// 	if (rst == 1'b1) begin
// 		dout <= 'b0 ;
// 	end
//     else begin
//     	for (m=0; m<32; m=m+1) begin 
//     		for (n=0; n<LUT_OUT_NUM_ONE_EQUATION; n=n+1) begin 
//     			if ( n<LUT_NUM_ONE_EQUATION ) begin
//     				dout[m*LUT_OUT_NUM_ONE_EQUATION+n] <= dout_pre[m*LUT_NUM_ONE_EQUATION+n];
//     			end
//     			else begin
//     				dout[m*LUT_OUT_NUM_ONE_EQUATION+n] <= 1'b0 ;
//     			end
//     		end
//     	end
//     end
// end

always @(posedge clk) begin

            dout <= dout_pre;

end

// always @(posedge clk) begin
//   if (rst == 1'b1) begin
//     dout <= 'b0 ;
//   end
//     else begin

//             dout <= dout_pre;
//           end

// end



endmodule 

// always @(posedge clk or posedge rst) begin
// 	if (rst == 1'b1) begin
// 		dout <= 'b0 ;
// 	end
//     else begin
//        dout <= dout_pre ; 
//     end
// end
// 
// parameter  [0:LUT_NUM_ONE_EQUATION*64*16-1] POLY  = { 
// 64'b1010101010101010101010101010101001010101010101011010101010101010,
// 64'b0011001100110011110011001100110001010101101010100101010110101010,
// 64'b0101101001011010010110100101101000001111111100000000111111110000,
// 64'b1100110011001100110011001100110000001111000011111111000011110000,
// 64'b1111111111111111000000000000000011000011110000110011110000111100,
// 64'b0110011010011001100110010110011000110011001100111100110011001100,
// 64'b0110100101101001100101101001011001011010010110100101101001011010,
// 64'b1111000011110000111100001111000001011010010110100101101001011010,
// 64'b1111111111111111000000000000000011111111111111110000000000000000,
// 64'b1010010101011010101001010101101011000011001111001100001100111100,
// 64'b1010101001010101010101011010101011001100110011001100110011001100,
// 64'b0101010110101010010101011010101000111100001111000011110000111100,
// 64'b1001100101100110100110010110011000000000000000000000000000000000,
// 64'b0110011001100110011001100110011011001100110011001100110011001100,
// 64'b1100001111000011001111000011110010011001100110010110011001100110,
// 64'b1100001100111100110000110011110000000000111111111111111100000000,
// 64'b0011110000111100001111000011110011111111000000001111111100000000,
// 64'b1111111111111111000000000000000010100101010110101010010101011010,
// 64'b0000111111110000000011111111000001011010010110100101101001011010,
// 64'b0000000011111111111111110000000010011001011001101001100101100110,
// 64'b1010010101011010101001010101101000110011110011000011001111001100,
// 64'b1111111111111111000000000000000000000000000000000000000000000000,
// 64'b1100001111000011001111000011110001011010101001011010010101011010,
// 64'b1001100101100110100110010110011011110000111100001111000011110000,
// 64'b1100110000110011001100111100110000001111111100000000111111110000,
// 64'b1010010101011010101001010101101000000000000000000000000000000000,
// 64'b1001011010010110100101101001011011110000111100001111000011110000,
// 64'b0011110011000011110000110011110000111100001111000011110000111100,
// 64'b0000000011111111111111110000000001010101010101011010101010101010,
// 64'b1100001100111100110000110011110001010101010101011010101010101010,
// 64'b1111111111111111000000000000000011001100001100110011001111001100,
// 64'b1100110011001100110011001100110000110011110011000011001111001100,
// 64'b1001011010010110100101101001011011000011110000110011110000111100,
// 64'b1001011001101001011010011001011000001111000011111111000011110000,
// 64'b1111111111111111000000000000000000000000000000000000000000000000,
// 64'b0000000000000000000000000000000011001100001100110011001111001100,
// 64'b1100001100111100110000110011110001010101101010100101010110101010,
// 64'b0101101010100101101001010101101000000000111111111111111100000000,
// 64'b0000000000000000000000000000000000000000000000000000000000000000,
// 64'b1100001100111100110000110011110011111111000000001111111100000000,
// 64'b1111000000001111000011111111000000001111111100000000111111110000,
// 64'b0101010101010101101010101010101011001100110011001100110011001100,
// 64'b0101101010100101101001010101101001100110011001100110011001100110,
// 64'b0000000000000000000000000000000010100101101001010101101001011010,
// 64'b0101101001011010010110100101101010100101101001010101101001011010,
// 64'b1100001100111100110000110011110000001111111100000000111111110000,
// 64'b0011110011000011110000110011110001010101101010100101010110101010,
// 64'b1010101010101010101010101010101010101010101010101010101010101010,
// 64'b1010101010101010101010101010101000001111000011111111000011110000,
// 64'b1111000000001111000011111111000010011001100110010110011001100110,
// 64'b1100110000110011001100111100110011111111111111110000000000000000,
// 64'b1010101010101010101010101010101010101010101010101010101010101010,
// 64'b0101101010100101101001010101101011111111111111110000000000000000,
// 64'b0011001111001100001100111100110000000000111111111111111100000000,
// 64'b0011110000111100001111000011110011110000111100001111000011110000,
// 64'b1010101001010101010101011010101000111100001111000011110000111100,
// 64'b0101010101010101101010101010101000110011110011000011001111001100,
// 64'b0101010101010101101010101010101010011001011001101001100101100110,
// 64'b1001100101100110100110010110011010101010010101010101010110101010,
// 64'b0000000011111111111111110000000000110011001100111100110011001100,
// 64'b1001100110011001011001100110011011001100110011001100110011001100,
// 64'b0110100110010110011010011001011011111111000000001111111100000000,
// 64'b1010101010101010101010101010101010010110100101101001011010010110,
// 64'b1111000000001111000011111111000010101010101010101010101010101010,
// 64'b1111111100000000111111110000000001100110011001100110011001100110,
// 64'b0110011010011001100110010110011000000000000000000000000000000000,
// 64'b1001011010010110100101101001011001010101010101011010101010101010,
// 64'b0101010110101010010101011010101001010101101010100101010110101010,
// 64'b1111111111111111000000000000000000001111111100000000111111110000,
// 64'b1001100110011001011001100110011000001111000011111111000011110000,
// 64'b0000000011111111111111110000000011000011110000110011110000111100,
// 64'b0000000000000000000000000000000000110011001100111100110011001100,
// 64'b0000111100001111111100001111000001011010010110100101101001011010,
// 64'b0110100101101001100101101001011001011010010110100101101001011010,
// 64'b0011001100110011110011001100110011111111111111110000000000000000,
// 64'b0110011010011001100110010110011011000011001111001100001100111100,
// 64'b0101010101010101101010101010101011001100110011001100110011001100,
// 64'b0011001111001100001100111100110000111100001111000011110000111100,
// 64'b1100001111000011001111000011110010101010101010101010101010101010,
// 64'b0110100110010110011010011001011011111111111111110000000000000000,
// 64'b0011001100110011110011001100110011000011110000110011110000111100,
// 64'b0000000000000000000000000000000011001100001100110011001111001100,
// 64'b1001011010010110100101101001011000000000111111111111111100000000,
// 64'b0101010101010101101010101010101011000011110000110011110000111100,
// 64'b1010101010101010101010101010101000110011001100111100110011001100,
// 64'b1111111100000000111111110000000001101001100101100110100110010110,
// 64'b0110100110010110011010011001011011001100001100110011001111001100,
// 64'b0101101001011010010110100101101010100101010110101010010101011010,
// 64'b0110100101101001100101101001011011110000111100001111000011110000,
// 64'b0110011001100110011001100110011010100101010110101010010101011010,
// 64'b0101101001011010010110100101101010010110100101101001011010010110,
// 64'b1010010101011010101001010101101001100110011001100110011001100110,
// 64'b1010010101011010101001010101101000110011001100111100110011001100,
// 64'b1010101010101010101010101010101011111111000000001111111100000000,
// 64'b0110011001100110011001100110011001101001011010011001011010010110,
// 64'b0011110011000011110000110011110010101010101010101010101010101010,
// 64'b1010101001010101010101011010101011000011110000110011110000111100,
// 64'b0000111100001111111100001111000000110011001100111100110011001100,
// 64'b0000111100001111111100001111000001100110100110011001100101100110,
// 64'b1100001100111100110000110011110011110000111100001111000011110000,
// 64'b1001011010010110100101101001011011000011110000110011110000111100,
// 64'b0110100101101001100101101001011001010101010101011010101010101010,
// 64'b1100001100111100110000110011110010011001100110010110011001100110,
// 64'b1010101010101010101010101010101001011010010110100101101001011010,
// 64'b0110011010011001100110010110011000111100001111000011110000111100,
// 64'b1111111100000000111111110000000011110000111100001111000011110000,
// 64'b1001011010010110100101101001011001010101010101011010101010101010,
// 64'b1111000011110000111100001111000011000011001111001100001100111100,
// 64'b0000111111110000000011111111000001100110011001100110011001100110,
// 64'b1111111100000000111111110000000000001111111100000000111111110000,
// 64'b0011110011000011110000110011110001011010010110100101101001011010,
// 64'b1010010101011010101001010101101001101001011010011001011010010110,
// 64'b1010010101011010101001010101101001010101101010100101010110101010,
// 64'b0110011001100110011001100110011000001111111100000000111111110000,
// 64'b0110100101101001100101101001011001100110011001100110011001100110,
// 64'b0000111100001111111100001111000010010110100101101001011010010110,
// 64'b0101010110101010010101011010101010011001011001101001100101100110,
// 64'b1100001111000011001111000011110000001111111100000000111111110000,
// 64'b0101010101010101101010101010101011111111000000001111111100000000,
// 64'b1100001100111100110000110011110011001100110011001100110011001100,
// 64'b1111111100000000111111110000000001011010101001011010010101011010,
// 64'b0000000011111111111111110000000000111100001111000011110000111100,
// 64'b1111111111111111000000000000000000000000111111111111111100000000,
// 64'b1111000000001111000011111111000000110011110011000011001111001100,
// 64'b0110011010011001100110010110011011000011001111001100001100111100,
// 64'b1100110000110011001100111100110010011001100110010110011001100110,
// 64'b0011110000111100001111000011110000000000111111111111111100000000,
// 64'b1100001100111100110000110011110000111100001111000011110000111100,
// 64'b0101010110101010010101011010101011000011001111001100001100111100,
// 64'b0110011001100110011001100110011000111100001111000011110000111100,
// 64'b1010010101011010101001010101101010101010010101010101010110101010,
// 64'b0101010101010101101010101010101011001100110011001100110011001100,
// 64'b0000000011111111111111110000000010101010101010101010101010101010,
// 64'b0011001100110011110011001100110000000000111111111111111100000000,
// 64'b0000000000000000000000000000000001011010101001011010010101011010,
// 64'b1100110000110011001100111100110010011001011001101001100101100110,
// 64'b1100001100111100110000110011110011001100110011001100110011001100,
// 64'b1001100110011001011001100110011000000000111111111111111100000000,
// 64'b0101101001011010010110100101101011000011110000110011110000111100,
// 64'b0000000000000000000000000000000011110000000011110000111111110000,
// 64'b0101101001011010010110100101101000001111000011111111000011110000,
// 64'b0110011010011001100110010110011010100101101001010101101001011010,
// 64'b1010010101011010101001010101101010010110100101101001011010010110,
// 64'b0110011010011001100110010110011000110011001100111100110011001100,
// 64'b1111111111111111000000000000000001011010010110100101101001011010,
// 64'b0000111100001111111100001111000011001100110011001100110011001100,
// 64'b1001011010010110100101101001011011111111111111110000000000000000,
// 64'b0101010101010101101010101010101001100110100110011001100101100110,
// 64'b0110100110010110011010011001011001101001011010011001011010010110,
// 64'b0011001111001100001100111100110011110000111100001111000011110000,
// 64'b1100110011001100110011001100110011111111111111110000000000000000,
// 64'b0110011010011001100110010110011010100101010110101010010101011010,
// 64'b1010010101011010101001010101101010101010010101010101010110101010,
// 64'b1001100110011001011001100110011001010101101010100101010110101010,
// 64'b1001011001101001011010011001011010011001011001101001100101100110,
// 64'b0000000000000000000000000000000001101001100101100110100110010110,
// 64'b0110100101101001100101101001011011110000111100001111000011110000,
// 64'b1001100110011001011001100110011010011001011001101001100101100110,
// 64'b0000111111110000000011111111000011110000111100001111000011110000,
// 64'b1010010101011010101001010101101000000000000000000000000000000000,
// 64'b0011001100110011110011001100110001101001011010011001011010010110,
// 64'b1111000011110000111100001111000001101001100101100110100110010110,
// 64'b0110011001100110011001100110011001010101101010100101010110101010,
// 64'b0000000000000000000000000000000000000000000000000000000000000000,
// 64'b0011110000111100001111000011110001100110100110011001100101100110,
// 64'b1100001111000011001111000011110000110011001100111100110011001100,
// 64'b1001011001101001011010011001011010011001100110010110011001100110,
// 64'b1100001111000011001111000011110011000011110000110011110000111100,
// 64'b0011001111001100001100111100110011000011001111001100001100111100,
// 64'b1100001100111100110000110011110011111111000000001111111100000000,
// 64'b1001011010010110100101101001011011000011110000110011110000111100,
// 64'b1010101001010101010101011010101011111111000000001111111100000000,
// 64'b1100110000110011001100111100110000000000000000000000000000000000,
// 64'b1111000011110000111100001111000011000011001111001100001100111100,
// 64'b0101010110101010010101011010101010010110011010010110100110010110,
// 64'b0011110000111100001111000011110000110011001100111100110011001100,
// 64'b0000000000000000000000000000000000000000000000000000000000000000,
// 64'b0000111111110000000011111111000011000011110000110011110000111100,
// 64'b0000111111110000000011111111000001011010010110100101101001011010,
// 64'b1001011001101001011010011001011010010110100101101001011010010110,
// 64'b1010010101011010101001010101101010100101010110101010010101011010,
// 64'b0101101001011010010110100101101010100101010110101010010101011010,
// 64'b1111000000001111000011111111000011111111111111110000000000000000,
// 64'b1100001100111100110000110011110000001111111100000000111111110000,
// 64'b0011001100110011110011001100110001010101010101011010101010101010,
// 64'b1010010110100101010110100101101000000000000000000000000000000000,
// 64'b0101010110101010010101011010101011110000000011110000111111110000,
// 64'b0011001100110011110011001100110000111100110000111100001100111100,
// 64'b0000111111110000000011111111000001011010010110100101101001011010,
// 64'b0000000000000000000000000000000010101010101010101010101010101010,
// 64'b0000000011111111111111110000000000001111111100000000111111110000,
// 64'b0000000011111111111111110000000010011001011001101001100101100110,
// 64'b0011110011000011110000110011110011000011001111001100001100111100,
// 64'b0110011010011001100110010110011011001100001100110011001111001100,
// 64'b0011001111001100001100111100110000110011110011000011001111001100,
// 64'b0000000011111111111111110000000000000000000000000000000000000000,
// 64'b0101101010100101101001010101101010101010010101010101010110101010,
// 64'b1111000011110000111100001111000011001100110011001100110011001100,
// 64'b1001100101100110100110010110011010101010101010101010101010101010,
// 64'b1001100110011001011001100110011000000000111111111111111100000000,
// 64'b1111000011110000111100001111000001011010101001011010010101011010,
// 64'b1010101001010101010101011010101010011001011001101001100101100110,
// 64'b0000000000000000000000000000000011001100110011001100110011001100,
// 64'b1111111111111111000000000000000000000000111111111111111100000000,
// 64'b0101010101010101101010101010101011000011110000110011110000111100,
// 64'b0101101010100101101001010101101011110000000011110000111111110000,
// 64'b0110100101101001100101101001011000001111000011111111000011110000,
// 64'b0101101001011010010110100101101001011010010110100101101001011010

//  } ; 