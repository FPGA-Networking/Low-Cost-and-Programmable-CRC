// **************************************************************
// COPYRIGHT(c)2015, Xidian University
// All rights reserved.
//
// IP LIB INDEX :  
// IP Name      :      
// File name    : 
// Module name  : 
// Full name    :  
//
// Author       : Liu-Huan 
// Email        : assasin9997@163.com 
// Data         : 
// Version      : V 1.0 
// 
// Abstract     : 
// Called by    :  
// 
// Modification history
// -----------------------------------------------------------------
// 
// 
//
// *****************************************************************

// *******************
// TIMESCALE
// ******************* 
`timescale 1ns/1ps 

// *******************
// INFORMATION
// *******************


//*******************
//DEFINE(s)
//*******************
//`define UDLY 1    //Unit delay, for non-blocking assignments in sequential logic



//*******************
//DEFINE MODULE PORT
//*******************
module  go_back_pipe 

# ( parameter   GO_BACK_STAGE        = 7      ,
                BUS_WIDTH            = 1024   ,
                MOD_WIDTH            = 7 

)

  (     
            input                       clk          ,
            input                       rst          ,
            input    [31:0]             crc_in       ,
            input                       crc_en_in    ,
            input    [MOD_WIDTH-1:0]    mod_in       ,
            output   [31:0]             crc_out      ,
            output                      crc_out_en
              ) ;

//*******************
//DEFINE LOCAL PARAMETER
//*******************
//parameter(s)
                                     
  parameter [0:GO_BACK_STAGE*32*64*6-1] POLY =                           
{
64'b1100110000110011110011000011001100110011110011000011001111001100,
64'b0011110000111100001111000011110000111100001111000011110000111100,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0110100110010110100101100110100110010110011010010110100110010110,
64'b1001100101100110100110010110011010011001011001101001100101100110,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1010010110100101010110100101101010100101101001010101101001011010,
64'b0101010101010101101010101010101001010101010101011010101010101010,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1100110000110011110011000011001100110011110011000011001111001100,
64'b0011001100110011001100110011001111001100110011001100110011001100,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1100001100111100001111001100001100111100110000111100001100111100,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0110100101101001100101101001011001101001011010011001011010010110,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0011110011000011001111001100001111000011001111001100001100111100,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b1111000011110000111100001111000011110000111100001111000011110000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1001011010010110011010010110100101101001011010011001011010010110,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b1111111100000000111111110000000011111111000000001111111100000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1111000011110000111100001111000011110000111100001111000011110000,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b1111111111111111000000000000000011111111111111110000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0101010110101010010101011010101001010101101010100101010110101010,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b1111111111111111111111111111111100000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0101010110101010101010100101010110101010010101010101010110101010,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000011111111111111110000000000000000111111111111111100000000,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1100110000110011001100111100110011001100001100110011001111001100,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1111000011110000111100001111000011110000111100001111000011110000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0101101001011010101001011010010110100101101001010101101001011010,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1111111100000000111111110000000011111111000000001111111100000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0110011010011001011001101001100110011001011001101001100101100110,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1111111111111111000000000000000011111111111111110000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0110100101101001100101101001011001101001011010011001011010010110,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1111111111111111111111111111111100000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0101101001011010010110100101101001011010010110100101101001011010,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1001100101100110100110010110011010011001011001101001100101100110,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1100001111000011001111000011110011000011110000110011110000111100,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1111000011110000111100001111000011110000111100001111000011110000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1111000000001111111100000000111100001111111100000000111111110000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1111111100000000111111110000000011111111000000001111111100000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1010101001010101010101011010101010101010010101010101010110101010,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1111111111111111000000000000000011111111111111110000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1100110011001100001100110011001100110011001100111100110011001100,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1111111111111111111111111111111100000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0110100110010110011010011001011001101001100101100110100110010110,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b0101101001011010101001011010010110100101101001010101101001011010,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b0110011010011001011001101001100110011001011001101001100101100110,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1100001111000011001111000011110011000011110000110011110000111100,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0011110000111100001111000011110000111100001111000011110000111100,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1010010101011010101001010101101010100101010110101010010101011010,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1100110000110011001100111100110011001100001100110011001111001100,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0101101001011010101001011010010110100101101001010101101001011010,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1100110000110011110011000011001100110011110011000011001111001100,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1010010110100101010110100101101010100101101001010101101001011010,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1010101010101010010101010101010101010101010101011010101010101010,
64'b1100110000110011110011000011001100110011110011000011001111001100,
64'b1100110000110011001100111100110011001100001100110011001111001100,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1001100110011001011001100110011010011001100110010110011001100110,
64'b0110100110010110100101100110100110010110011010010110100110010110,
64'b1001011001101001100101100110100101101001100101100110100110010110,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1100001111000011001111000011110011000011110000110011110000111100,
64'b0000111100001111111100001111000000001111000011111111000011110000,
64'b0101101001011010010110100101101001011010010110100101101001011010,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0101101010100101010110101010010110100101010110101010010101011010,
64'b0000000011111111000000001111111111111111000000001111111100000000,
64'b0011001111001100001100111100110000110011110011000011001111001100,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1100110000110011110011000011001100110011110011000011001111001100,
64'b1001100101100110011001101001100101100110100110011001100101100110,
64'b0110100110010110011010011001011001101001100101100110100110010110,
64'b1111000011110000111100001111000011110000111100001111000011110000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1010010110100101101001011010010101011010010110100101101001011010,
64'b0101101010100101101001010101101001011010101001011010010101011010,
64'b0101101001011010010110100101101001011010010110100101101001011010,
64'b1111111100000000111111110000000011111111000000001111111100000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1001100101100110100110010110011010011001011001101001100101100110,
64'b1001100101100110011001101001100101100110100110011001100101100110,
64'b0011001111001100001100111100110000110011110011000011001111001100,
64'b1111111111111111000000000000000011111111111111110000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0110100101101001011010010110100110010110100101101001011010010110,
64'b1111000000001111000011111111000011110000000011110000111111110000,
64'b0110100110010110011010011001011001101001100101100110100110010110,
64'b1111111111111111111111111111111100000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1100001100111100001111001100001100111100110000111100001100111100,
64'b1001100110011001011001100110011010011001100110010110011001100110,
64'b1111000011110000111100001111000011110000111100001111000011110000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000111111110000111100000000111111110000000011110000111111110000,
64'b0110100101101001011010010110100110010110100101101001011010010110,
64'b1111111100000000111111110000000011111111000000001111111100000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1111111100000000111111110000000011111111000000001111111100000000,
64'b1010010110100101101001011010010101011010010110100101101001011010,
64'b1001100101100110100110010110011010011001011001101001100101100110,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1111000011110000111100001111000011110000111100001111000011110000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0101010101010101010101010101010110101010101010101010101010101010,
64'b1111111111111111111111111111111100000000000000000000000000000000,
64'b1010010101011010101001010101101010100101010110101010010101011010,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1111111100000000111111110000000011111111000000001111111100000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1100110011001100001100110011001100110011001100111100110011001100,
64'b0110011010011001011001101001100110011001011001101001100101100110,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1111111111111111000000000000000011111111111111110000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000111100001111000011110000111111110000111100001111000011110000,
64'b0110100101101001100101101001011001101001011010011001011010010110,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1111111111111111111111111111111100000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0101010110101010010101011010101001010101101010100101010110101010,
64'b1001011001101001100101100110100101101001100101100110100110010110,
64'b0011110000111100001111000011110000111100001111000011110000111100,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b0011001100110011110011001100110000110011001100111100110011001100,
64'b0011110011000011110000110011110000111100110000111100001100111100,
64'b1010010101011010101001010101101010100101010110101010010101011010,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b0000111100001111111100001111000000001111000011111111000011110000,
64'b1100001111000011001111000011110011000011110000110011110000111100,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1010101001010101101010100101010101010101101010100101010110101010,
64'b1111000000001111111100000000111100001111111100000000111111110000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0011001100110011110011001100110000110011001100111100110011001100,
64'b1010101001010101010101011010101010101010010101010101010110101010,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1010010110100101101001011010010101011010010110100101101001011010,
64'b1100110011001100001100110011001100110011001100111100110011001100,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0011001111001100001100111100110000110011110011000011001111001100,
64'b1010010110100101101001011010010101011010010110100101101001011010,
64'b0101101001011010010110100101101001011010010110100101101001011010,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000111100001111111100001111000000001111000011111111000011110000,
64'b0011001111001100001100111100110000110011110011000011001111001100,
64'b1001100101100110100110010110011010011001011001101001100101100110,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1010101001010101010101011010101010101010010101010101010110101010,
64'b1100001100111100001111001100001100111100110000111100001100111100,
64'b0000111111110000000011111111000000001111111100000000111111110000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b1100001111000011001111000011110011000011110000110011110000111100,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0011110000111100001111000011110000111100001111000011110000111100,
64'b1111000000001111111100000000111100001111111100000000111111110000,
64'b0011110000111100001111000011110000111100001111000011110000111100,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1010010101011010101001010101101010100101010110101010010101011010,
64'b0000000011111111111111110000000000000000111111111111111100000000,
64'b1010010101011010101001010101101010100101010110101010010101011010,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1100110000110011110011000011001100110011110011000011001111001100,
64'b1100110000110011001100111100110011001100001100110011001111001100,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1010010110100101010110100101101010100101101001010101101001011010,
64'b0101101001011010101001011010010110100101101001010101101001011010,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0110011010011001011001101001100110011001011001101001100101100110,
64'b1100110000110011110011000011001100110011110011000011001111001100,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1100001111000011001111000011110011000011110000110011110000111100,
64'b1010010110100101010110100101101010100101101001010101101001011010,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1111000000001111111100000000111100001111111100000000111111110000,
64'b1100110000110011110011000011001100110011110011000011001111001100,
64'b0011110000111100001111000011110000111100001111000011110000111100,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000011111111111111110000000000000000111111111111111100000000,
64'b1010010110100101010110100101101010100101101001010101101001011010,
64'b1010010101011010101001010101101010100101010110101010010101011010,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1100001111000011110000111100001100111100001111000011110000111100,
64'b1111111100000000111111110000000011111111000000001111111100000000,
64'b0000111100001111111100001111000000001111000011111111000011110000,
64'b1111000000001111111100000000111100001111111100000000111111110000,
64'b1100110000110011110011000011001100110011110011000011001111001100,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b0110011010011001011001101001100110011001011001101001100101100110,
64'b1010101001010101010101011010101010101010010101010101010110101010,
64'b0000111111110000111100000000111111110000000011110000111111110000,
64'b1111000011110000000011110000111100001111000011111111000011110000,
64'b0110100110010110100101100110100110010110011010010110100110010110,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b0000000000000000111111111111111111111111111111110000000000000000,
64'b1001100101100110011001101001100101100110100110011001100101100110,
64'b1111000000001111111100000000111100001111111100000000111111110000,
64'b0101101001011010010110100101101001011010010110100101101001011010,
64'b1010010110100101010110100101101010100101101001010101101001011010,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b0101010101010101010101010101010110101010101010101010101010101010,
64'b1001011010010110011010010110100101101001011010011001011010010110,
64'b1010101001010101010101011010101010101010010101010101010110101010,
64'b1001100101100110100110010110011010011001011001101001100101100110,
64'b1100110000110011110011000011001100110011110011000011001111001100,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b1010010110100101101001011010010101011010010110100101101001011010,
64'b0110100101101001011010010110100110010110100101101001011010010110,
64'b0110100101101001011010010110100110010110100101101001011010010110,
64'b0011001111001100110011000011001111001100001100110011001111001100,
64'b1100001100111100001111001100001100111100110000111100001100111100,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b1111000000001111111100000000111100001111111100000000111111110000,
64'b1001011010010110100101101001011010010110100101101001011010010110,
64'b0110011010011001100110010110011001100110100110011001100101100110,
64'b1010101001010101010101011010101010101010010101010101010110101010,
64'b0110100101101001100101101001011001101001011010011001011010010110,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b1010101001010101010101011010101010101010010101010101010110101010,
64'b0110100110010110011010011001011001101001100101100110100110010110,
64'b0011110000111100110000111100001111000011110000110011110000111100,
64'b1100110011001100001100110011001100110011001100111100110011001100,
64'b0011110011000011001111001100001111000011001111001100001100111100,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b1010010110100101010110100101101010100101101001010101101001011010,
64'b1100001111000011001111000011110011000011110000110011110000111100,
64'b1111111100000000000000001111111100000000111111111111111100000000,
64'b0101010110101010010101011010101001010101101010100101010110101010,
64'b1001011010010110011010010110100101101001011010011001011010010110,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b0000111111110000000011111111000000001111111100000000111111110000,
64'b0000111100001111000011110000111111110000111100001111000011110000,
64'b0000111100001111000011110000111111110000111100001111000011110000,
64'b0110100110010110100101100110100110010110011010010110100110010110,
64'b1111000011110000111100001111000011110000111100001111000011110000,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b0000000011111111111111110000000000000000111111111111111100000000,
64'b1111111100000000111111110000000011111111000000001111111100000000,
64'b0101010110101010010101011010101001010101101010100101010110101010,
64'b0110100110010110100101100110100110010110011010010110100110010110,
64'b0101010110101010010101011010101001010101101010100101010110101010,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b0110100101101001100101101001011001101001011010011001011010010110,
64'b0000000011111111111111110000000000000000111111111111111100000000,
64'b0011110000111100001111000011110000111100001111000011110000111100,
64'b0011001100110011110011001100110000110011001100111100110011001100,
64'b0101010110101010101010100101010110101010010101010101010110101010,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b0101010110101010010101011010101001010101101010100101010110101010,
64'b1111111100000000000000001111111100000000111111111111111100000000,
64'b0000000011111111111111110000000000000000111111111111111100000000,
64'b1111111100000000111111110000000011111111000000001111111100000000,
64'b0000000011111111111111110000000000000000111111111111111100000000,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b1111000011110000000011110000111100001111000011111111000011110000,
64'b1111111100000000000000001111111100000000111111111111111100000000,
64'b1010010110100101101001011010010101011010010110100101101001011010,
64'b0000111111110000111100000000111111110000000011110000111111110000,
64'b1100110000110011001100111100110011001100001100110011001111001100,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1010101001010101101010100101010101010101101010100101010110101010,
64'b1010101010101010010101010101010101010101010101011010101010101010,
64'b1001100101100110100110010110011010011001011001101001100101100110,
64'b0101010110101010101010100101010110101010010101010101010110101010,
64'b0101101001011010101001011010010110100101101001010101101001011010,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0011001100110011110011001100110000110011001100111100110011001100,
64'b1001100110011001100110011001100101100110011001100110011001100110,
64'b0110100101101001100101101001011001101001011010011001011010010110,
64'b1100110011001100001100110011001100110011001100111100110011001100,
64'b0110011010011001011001101001100110011001011001101001100101100110,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b1010010110100101101001011010010101011010010110100101101001011010,
64'b0011110000111100001111000011110000111100001111000011110000111100,
64'b1001011001101001100101100110100101101001100101100110100110010110,
64'b0000111100001111000011110000111111110000111100001111000011110000,
64'b0110100101101001100101101001011001101001011010011001011010010110,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b0101101010100101010110101010010110100101010110101010010101011010,
64'b0101101001011010010110100101101001011010010110100101101001011010,
64'b0011001111001100001100111100110000110011110011000011001111001100,
64'b1010010110100101101001011010010101011010010110100101101001011010,
64'b0101101001011010010110100101101001011010010110100101101001011010,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1100110000110011001100111100110011001100001100110011001111001100,
64'b1001100101100110100110010110011010011001011001101001100101100110,
64'b0000111100001111111100001111000000001111000011111111000011110000,
64'b0011001111001100001100111100110000110011110011000011001111001100,
64'b1001100101100110100110010110011010011001011001101001100101100110,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1111000011110000000011110000111100001111000011111111000011110000,
64'b1100001111000011001111000011110011000011110000110011110000111100,
64'b0000000011111111000000001111111111111111000000001111111100000000,
64'b0000111100001111111100001111000000001111000011111111000011110000,
64'b1100001111000011001111000011110011000011110000110011110000111100,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000011111111000000001111111111111111000000001111111100000000,
64'b0101101010100101010110101010010110100101010110101010010101011010,
64'b1111111111111111000000000000000011111111111111110000000000000000,
64'b1010101001010101101010100101010101010101101010100101010110101010,
64'b1111000000001111111100000000111100001111111100000000111111110000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0101010101010101101010101010101001010101010101011010101010101010,
64'b0110011010011001100110010110011001100110100110011001100101100110,
64'b0101010101010101010101010101010110101010101010101010101010101010,
64'b0011001100110011110011001100110000110011001100111100110011001100,
64'b1010101001010101010101011010101010101010010101010101010110101010,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b1001100110011001100110011001100101100110011001100110011001100110,
64'b0011110000111100110000111100001111000011110000110011110000111100,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b1010010110100101101001011010010101011010010110100101101001011010,
64'b1100110011001100001100110011001100110011001100111100110011001100,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b0101010101010101010101010101010110101010101010101010101010101010,
64'b1010010110100101101001011010010101011010010110100101101001011010,
64'b0101010101010101101010101010101001010101010101011010101010101010,
64'b1100001111000011110000111100001100111100001111000011110000111100,
64'b0110100110010110011010011001011001101001100101100110100110010110,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b1010010110100101101001011010010101011010010110100101101001011010,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b1001011010010110011010010110100101101001011010011001011010010110,
64'b1111111111111111111111111111111100000000000000000000000000000000,
64'b0101101001011010101001011010010110100101101001010101101001011010,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1001100101100110100110010110011010011001011001101001100101100110,
64'b1001011010010110100101101001011010010110100101101001011010010110,
64'b0011110011000011001111001100001111000011001111001100001100111100,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b0110011010011001011001101001100110011001011001101001100101100110,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b0110100101101001100101101001011001101001011010011001011010010110,
64'b1100001100111100110000110011110011000011001111001100001100111100,
64'b1111000000001111000011111111000011110000000011110000111111110000,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b1100001111000011001111000011110011000011110000110011110000111100,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b1111111100000000111111110000000011111111000000001111111100000000,
64'b0000111100001111111100001111000000001111000011111111000011110000,
64'b1111000000001111111100000000111100001111111100000000111111110000,
64'b1100110000110011110011000011001100110011110011000011001111001100,
64'b0011110000111100001111000011110000111100001111000011110000111100,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0101010101010101101010101010101001010101010101011010101010101010,
64'b0000000011111111000000001111111111111111000000001111111100000000,
64'b0000000011111111111111110000000000000000111111111111111100000000,
64'b1010010110100101010110100101101010100101101001010101101001011010,
64'b1010010101011010101001010101101010100101010110101010010101011010,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0011001100110011001100110011001111001100110011001100110011001100,
64'b1111111111111111000000000000000011111111111111110000000000000000,
64'b1010101010101010010101010101010101010101010101011010101010101010,
64'b1100110000110011110011000011001100110011110011000011001111001100,
64'b1100110000110011001100111100110011001100001100110011001111001100,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1111000011110000111100001111000011110000111100001111000011110000,
64'b0101010101010101010101010101010110101010101010101010101010101010,
64'b0011001100110011001100110011001111001100110011001100110011001100,
64'b1010010110100101010110100101101010100101101001010101101001011010,
64'b0101101001011010101001011010010110100101101001010101101001011010,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0101010110101010010101011010101001010101101010100101010110101010,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b0101101001011010010110100101101001011010010110100101101001011010,
64'b0110011010011001011001101001100110011001011001101001100101100110,
64'b1100110000110011110011000011001100110011110011000011001111001100,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b1001100110011001011001100110011010011001100110010110011001100110,
64'b1111000011110000111100001111000011110000111100001111000011110000,
64'b0011001111001100001100111100110000110011110011000011001111001100,
64'b1100001111000011001111000011110011000011110000110011110000111100,
64'b1010010110100101010110100101101010100101101001010101101001011010,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b1100001111000011001111000011110011000011110000110011110000111100,
64'b1100001111000011110000111100001100111100001111000011110000111100,
64'b0110100101101001011010010110100110010110100101101001011010010110,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b0110100110010110100101100110100110010110011010010110100110010110,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b0011001111001100110011000011001111001100001100110011001111001100,
64'b1100110000110011110011000011001100110011110011000011001111001100,
64'b0000000011111111000000001111111111111111000000001111111100000000,
64'b1001011010010110100101101001011010010110100101101001011010010110,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1001100110011001100110011001100101100110011001100110011001100110,
64'b0110011001100110100110011001100110011001100110010110011001100110,
64'b0011110000111100110000111100001111000011110000110011110000111100,
64'b1010010101011010101001010101101010100101010110101010010101011010,
64'b1010010101011010010110101010010101011010101001011010010101011010,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b0011110000111100001111000011110000111100001111000011110000111100,
64'b0110100101101001011010010110100110010110100101101001011010010110,
64'b0101101010100101010110101010010110100101010110101010010101011010,
64'b0110011010011001100110010110011001100110100110011001100101100110,
64'b0011001111001100110011000011001111001100001100110011001111001100,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b0110011010011001100110010110011001100110100110011001100101100110,
64'b0000000011111111000000001111111111111111000000001111111100000000,
64'b0000111111110000111100000000111111110000000011110000111111110000,
64'b0101101001011010101001011010010110100101101001010101101001011010,
64'b1001100101100110100110010110011010011001011001101001100101100110,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0101010101010101010101010101010110101010101010101010101010101010,
64'b0011110000111100110000111100001111000011110000110011110000111100,
64'b0011110011000011110000110011110000111100110000111100001100111100,
64'b1010101001010101101010100101010101010101101010100101010110101010,
64'b0000000011111111000000001111111111111111000000001111111100000000,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b0101101010100101010110101010010110100101010110101010010101011010,
64'b1010010101011010010110101010010101011010101001011010010101011010,
64'b0011001100110011110011001100110000110011001100111100110011001100,
64'b0101010101010101101010101010101001010101010101011010101010101010,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b1111111111111111000000000000000011111111111111110000000000000000,
64'b0000111111110000111100000000111111110000000011110000111111110000,
64'b1111000000001111000011111111000011110000000011110000111111110000,
64'b0110100101101001011010010110100110010110100101101001011010010110,
64'b0101101010100101101001010101101001011010101001011010010101011010,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b1001011010010110011010010110100101101001011010011001011010010110,
64'b0011110011000011110000110011110000111100110000111100001100111100,
64'b0011110011000011110000110011110000111100110000111100001100111100,
64'b0000111111110000000011111111000000001111111100000000111111110000,
64'b1111000011110000111100001111000011110000111100001111000011110000,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b0011110011000011001111001100001111000011001111001100001100111100,
64'b1010010101011010010110101010010101011010101001011010010101011010,
64'b0000111111110000111100000000111111110000000011110000111111110000,
64'b0000000011111111111111110000000000000000111111111111111100000000,
64'b1111111100000000111111110000000011111111000000001111111100000000,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b0011001111001100001100111100110000110011110011000011001111001100,
64'b0101101010100101101001010101101001011010101001011010010101011010,
64'b0011110011000011110000110011110000111100110000111100001100111100,
64'b0110011001100110100110011001100110011001100110010110011001100110,
64'b1001011001101001100101100110100101101001100101100110100110010110,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b1111000000001111000011111111000011110000000011110000111111110000,
64'b0110011010011001100110010110011001100110100110011001100101100110,
64'b0000111100001111000011110000111111110000111100001111000011110000,
64'b1111111111111111111111111111111100000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0101010101010101101010101010101001010101010101011010101010101010,
64'b0011110011000011110000110011110000111100110000111100001100111100,
64'b0101010101010101101010101010101001010101010101011010101010101010,
64'b0011001111001100001100111100110000110011110011000011001111001100,
64'b1100001100111100001111001100001100111100110000111100001100111100,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b0011001100110011001100110011001111001100110011001100110011001100,
64'b0000111111110000111100000000111111110000000011110000111111110000,
64'b0011001100110011001100110011001111001100110011001100110011001100,
64'b0000111100001111111100001111000000001111000011111111000011110000,
64'b0000111111110000111100000000111111110000000011110000111111110000,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b0101101001011010010110100101101001011010010110100101101001011010,
64'b0101010110101010101010100101010110101010010101010101010110101010,
64'b0101101001011010010110100101101001011010010110100101101001011010,
64'b1010101001010101101010100101010101010101101010100101010110101010,
64'b1111111100000000000000001111111100000000111111111111111100000000,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b1001100101100110100110010110011010011001011001101001100101100110,
64'b1100110011001100001100110011001100110011001100111100110011001100,
64'b1001100101100110100110010110011010011001011001101001100101100110,
64'b0011001100110011110011001100110000110011001100111100110011001100,
64'b1010101010101010010101010101010101010101010101011010101010101010,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b0000000000000000111111111111111111111111111111110000000000000000,
64'b1100001111000011110000111100001100111100001111000011110000111100,
64'b0101101010100101101001010101101001011010101001011010010101011010,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b1111000011110000111100001111000011110000111100001111000011110000,
64'b1111111111111111111111111111111100000000000000000000000000000000,
64'b1010010101011010101001010101101010100101010110101010010101011010,
64'b1001100101100110011001101001100101100110100110011001100101100110,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0101101001011010010110100101101001011010010110100101101001011010,
64'b1111111100000000111111110000000011111111000000001111111100000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0110011010011001100110010110011001100110100110011001100101100110,
64'b0011110000111100110000111100001111000011110000110011110000111100,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b1001100101100110100110010110011010011001011001101001100101100110,
64'b1111111111111111000000000000000011111111111111110000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0011110000111100110000111100001111000011110000110011110000111100,
64'b1111000000001111111100000000111100001111111100000000111111110000,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b1100001111000011001111000011110011000011110000110011110000111100,
64'b1111111111111111111111111111111100000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1111000000001111111100000000111100001111111100000000111111110000,
64'b1010101001010101010101011010101010101010010101010101010110101010,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b0101101010100101010110101010010110100101010110101010010101011010,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b0000000011111111111111110000000000000000111111111111111100000000,
64'b0110011001100110100110011001100110011001100110010110011001100110,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b0000111111110000000011111111000000001111111100000000111111110000,
64'b0110100101101001011010010110100110010110100101101001011010010110,
64'b1010010110100101101001011010010101011010010110100101101001011010,
64'b1100110011001100001100110011001100110011001100111100110011001100,
64'b1010101001010101010101011010101010101010010101010101010110101010,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b1100001100111100110000110011110011000011001111001100001100111100,
64'b0000000011111111000000001111111111111111000000001111111100000000,
64'b1111000000001111111100000000111100001111111100000000111111110000,
64'b0110100101101001011010010110100110010110100101101001011010010110,
64'b0000111111110000000011111111000000001111111100000000111111110000,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b1111000000001111000011111111000011110000000011110000111111110000,
64'b1111111111111111000000000000000011111111111111110000000000000000,
64'b1010101001010101010101011010101010101010010101010101010110101010,
64'b0110100110010110011010011001011001101001100101100110100110010110,
64'b1010101001010101010101011010101010101010010101010101010110101010,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b1111111100000000000000001111111100000000111111111111111100000000,
64'b1111111111111111111111111111111100000000000000000000000000000000,
64'b1100110011001100001100110011001100110011001100111100110011001100,
64'b0011110011000011110000110011110000111100110000111100001100111100,
64'b1100110011001100001100110011001100110011001100111100110011001100,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1100001111000011110000111100001100111100001111000011110000111100,
64'b0110100101101001011010010110100110010110100101101001011010010110,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b0110100110010110100101100110100110010110011010010110100110010110,
64'b0110011010011001100110010110011001100110100110011001100101100110,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b0000111111110000000011111111000000001111111100000000111111110000,
64'b0110100110010110011010011001011001101001100101100110100110010110,
64'b0101101001011010010110100101101001011010010110100101101001011010,
64'b1100001100111100001111001100001100111100110000111100001100111100,
64'b1001011010010110011010010110100101101001011010011001011010010110,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1010101001010101010101011010101010101010010101010101010110101010,
64'b0011110011000011110000110011110000111100110000111100001100111100,
64'b0011001111001100001100111100110000110011110011000011001111001100,
64'b0000111111110000111100000000111111110000000011110000111111110000,
64'b1001011001101001100101100110100101101001100101100110100110010110,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b1100110011001100001100110011001100110011001100111100110011001100,
64'b0000111111110000111100000000111111110000000011110000111111110000,
64'b0000111100001111111100001111000000001111000011111111000011110000,
64'b1111111100000000000000001111111100000000111111111111111100000000,
64'b1001011001101001011010011001011010010110011010010110100110010110,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b1010010110100101101001011010010101011010010110100101101001011010,
64'b0101010110101010101010100101010110101010010101010101010110101010,
64'b1010101001010101101010100101010101010101101010100101010110101010,
64'b0000000000000000111111111111111111111111111111110000000000000000,
64'b0110100110010110100101100110100110010110011010010110100110010110,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b1001100101100110100110010110011010011001011001101001100101100110,
64'b0110011001100110100110011001100110011001100110010110011001100110,
64'b1001100110011001011001100110011010011001100110010110011001100110,
64'b0101010101010101010101010101010110101010101010101010101010101010,
64'b0110100110010110100101100110100110010110011010010110100110010110,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b0011001100110011110011001100110000110011001100111100110011001100,
64'b0000000000000000111111111111111111111111111111110000000000000000,
64'b1010010110100101101001011010010101011010010110100101101001011010,
64'b0101010110101010101010100101010110101010010101010101010110101010,
64'b0000111100001111111100001111000000001111000011111111000011110000,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b0011110000111100110000111100001111000011110000110011110000111100,
64'b1111111111111111000000000000000011111111111111110000000000000000,
64'b0011110011000011001111001100001111000011001111001100001100111100,
64'b0011001111001100001100111100110000110011110011000011001111001100,
64'b1010010101011010010110101010010101011010101001011010010101011010,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b1100001100111100001111001100001100111100110000111100001100111100,
64'b0101010101010101101010101010101001010101010101011010101010101010,
64'b0101010110101010101010100101010110101010010101010101010110101010,
64'b1111000000001111111100000000111100001111111100000000111111110000,
64'b0011110011000011001111001100001111000011001111001100001100111100,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b1010010101011010010110101010010101011010101001011010010101011010,
64'b1001100110011001100110011001100101100110011001100110011001100110,
64'b1100110011001100001100110011001100110011001100111100110011001100,
64'b1010101001010101010101011010101010101010010101010101010110101010,
64'b0101101010100101101001010101101001011010101001011010010101011010,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b0000000011111111000000001111111111111111000000001111111100000000,
64'b1001011010010110011010010110100101101001011010011001011010010110,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0011001111001100001100111100110000110011110011000011001111001100,
64'b0011110011000011001111001100001111000011001111001100001100111100,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b1001011001101001011010011001011010010110011010010110100110010110,
64'b0000111100001111000011110000111111110000111100001111000011110000,
64'b0101101010100101010110101010010110100101010110101010010101011010,
64'b1111111100000000111111110000000011111111000000001111111100000000,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b0101101001011010010110100101101001011010010110100101101001011010,
64'b1100001100111100001111001100001100111100110000111100001100111100,
64'b1111111100000000111111110000000011111111000000001111111100000000,
64'b0110011010011001100110010110011001100110100110011001100101100110,
64'b0101010101010101101010101010101001010101010101011010101010101010,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000011111111111111110000000000000000111111111111111100000000,
64'b0000111111110000000011111111000000001111111100000000111111110000,
64'b1111000011110000000011110000111100001111000011111111000011110000,
64'b0110100110010110011010011001011001101001100101100110100110010110,
64'b0011110000111100110000111100001111000011110000110011110000111100,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b1001100110011001100110011001100101100110011001100110011001100110,
64'b0000000011111111000000001111111111111111000000001111111100000000,
64'b1010010101011010101001010101101010100101010110101010010101011010,
64'b1100001111000011110000111100001100111100001111000011110000111100,
64'b1111111100000000000000001111111100000000111111111111111100000000,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b0011110000111100001111000011110000111100001111000011110000111100,
64'b0101010101010101101010101010101001010101010101011010101010101010,
64'b0110011010011001100110010110011001100110100110011001100101100110,
64'b0000111111110000000011111111000000001111111100000000111111110000,
64'b1010101010101010010101010101010101010101010101011010101010101010,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b1001011001101001011010011001011010010110011010010110100110010110,
64'b0011001100110011110011001100110000110011001100111100110011001100,
64'b1001100110011001011001100110011010011001100110010110011001100110,
64'b0101010101010101010101010101010110101010101010101010101010101010,
64'b0011110000111100110000111100001111000011110000110011110000111100,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b1111000000001111111100000000111100001111111100000000111111110000,
64'b0000111100001111111100001111000000001111000011111111000011110000,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b1001100101100110011001101001100101100110100110011001100101100110,
64'b0101010110101010101010100101010110101010010101010101010110101010,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0011001111001100001100111100110000110011110011000011001111001100,
64'b1010101001010101010101011010101010101010010101010101010110101010,
64'b1001100110011001100110011001100101100110011001100110011001100110,
64'b0110100110010110011010011001011001101001100101100110100110010110,
64'b0110100101101001011010010110100110010110100101101001011010010110,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1010010110100101010110100101101010100101101001010101101001011010,
64'b1100110011001100001100110011001100110011001100111100110011001100,
64'b0011110000111100001111000011110000111100001111000011110000111100,
64'b1001011001101001011010011001011010010110011010010110100110010110,
64'b1100001100111100110000110011110011000011001111001100001100111100,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b1100110000110011110011000011001100110011110011000011001111001100,
64'b0000111100001111000011110000111111110000111100001111000011110000,
64'b1010010101011010101001010101101010100101010110101010010101011010,
64'b1100001100111100001111001100001100111100110000111100001100111100,
64'b1111000000001111000011111111000011110000000011110000111111110000,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b1010010110100101010110100101101010100101101001010101101001011010,
64'b0101010110101010010101011010101001010101101010100101010110101010,
64'b0110011010011001100110010110011001100110100110011001100101100110,
64'b0000111111110000111100000000111111110000000011110000111111110000,
64'b0101010110101010101010100101010110101010010101010101010110101010,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0101010110101010101010100101010110101010010101010101010110101010,
64'b0011001100110011001100110011001111001100110011001100110011001100,
64'b1001100110011001011001100110011010011001100110010110011001100110,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b0110100101101001011010010110100110010110100101101001011010010110,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1100110011001100001100110011001100110011001100111100110011001100,
64'b0101101001011010010110100101101001011010010110100101101001011010,
64'b0110100101101001011010010110100110010110100101101001011010010110,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b1100001100111100110000110011110011000011001111001100001100111100,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b0000111100001111000011110000111111110000111100001111000011110000,
64'b1001100101100110100110010110011010011001011001101001100101100110,
64'b1100001100111100110000110011110011000011001111001100001100111100,
64'b0101101001011010010110100101101001011010010110100101101001011010,
64'b1111000000001111000011111111000011110000000011110000111111110000,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b0101010110101010010101011010101001010101101010100101010110101010,
64'b0110100101101001100101101001011001101001011010011001011010010110,
64'b1111000000001111000011111111000011110000000011110000111111110000,
64'b0011001111001100001100111100110000110011110011000011001111001100,
64'b1111111100000000000000001111111100000000111111111111111100000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1001100110011001011001100110011010011001100110010110011001100110,
64'b0011110011000011001111001100001111000011001111001100001100111100,
64'b1111111100000000000000001111111100000000111111111111111100000000,
64'b0000111100001111111100001111000000001111000011111111000011110000,
64'b0000000000000000111111111111111111111111111111110000000000000000,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b1100001111000011110000111100001100111100001111000011110000111100,
64'b1111000000001111000011111111000011110000000011110000111111110000,
64'b1010101010101010010101010101010101010101010101011010101010101010,
64'b1010101001010101101010100101010101010101101010100101010110101010,
64'b1111111111111111111111111111111100000000000000000000000000000000,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b1001011001101001011010011001011010010110011010010110100110010110,
64'b0101010110101010010101011010101001010101101010100101010110101010,
64'b1001011010010110100101101001011010010110100101101001011010010110,
64'b1100110000110011110011000011001100110011110011000011001111001100,
64'b1010010110100101010110100101101010100101101001010101101001011010,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b1111000000001111111100000000111100001111111100000000111111110000,
64'b0011001100110011001100110011001111001100110011001100110011001100,
64'b0110011010011001011001101001100110011001011001101001100101100110,
64'b0101101010100101010110101010010110100101010110101010010101011010,
64'b0110100110010110100101100110100110010110011010010110100110010110,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b0000000011111111111111110000000000000000111111111111111100000000,
64'b0101101001011010010110100101101001011010010110100101101001011010,
64'b0110100101101001100101101001011001101001011010011001011010010110,
64'b0110011010011001100110010110011001100110100110011001100101100110,
64'b0110100110010110100101100110100110010110011010010110100110010110,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b1010101010101010010101010101010101010101010101011010101010101010,
64'b0011001111001100001100111100110000110011110011000011001111001100,
64'b0011110011000011001111001100001111000011001111001100001100111100,
64'b0011110000111100110000111100001111000011110000110011110000111100,
64'b1100001100111100001111001100001100111100110000111100001100111100,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b0000000000000000111111111111111111111111111111110000000000000000,
64'b1010010110100101101001011010010101011010010110100101101001011010,
64'b0101010110101010101010100101010110101010010101010101010110101010,
64'b0000111100001111111100001111000000001111000011111111000011110000,
64'b1010101001010101101010100101010101010101101010100101010110101010,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b1111111111111111111111111111111100000000000000000000000000000000,
64'b1001100101100110100110010110011010011001011001101001100101100110,
64'b0110011001100110100110011001100110011001100110010110011001100110,
64'b1010101001010101101010100101010101010101101010100101010110101010,
64'b0011001100110011110011001100110000110011001100111100110011001100,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b0110100101101001100101101001011001101001011010011001011010010110,
64'b1100001111000011110000111100001100111100001111000011110000111100,
64'b1001100110011001011001100110011010011001100110010110011001100110,
64'b1010010110100101101001011010010101011010010110100101101001011010,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b0011110011000011001111001100001111000011001111001100001100111100,
64'b0000111111110000000011111111000000001111111100000000111111110000,
64'b0110100101101001011010010110100110010110100101101001011010010110,
64'b0011001111001100001100111100110000110011110011000011001111001100,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b1111000011110000111100001111000011110000111100001111000011110000,
64'b1111000000001111000011111111000011110000000011110000111111110000,
64'b1010101001010101010101011010101010101010010101010101010110101010,
64'b1100001100111100110000110011110011000011001111001100001100111100,
64'b1010010110100101010110100101101010100101101001010101101001011010,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b0101010110101010010101011010101001010101101010100101010110101010,
64'b1111111100000000000000001111111100000000111111111111111100000000,
64'b1100110011001100001100110011001100110011001100111100110011001100,
64'b1111000000001111000011111111000011110000000011110000111111110000,
64'b1100110000110011110011000011001100110011110011000011001111001100,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1001100101100110011001101001100101100110100110011001100101100110,
64'b1001100101100110100110010110011010011001011001101001100101100110,
64'b0011001100110011001100110011001111001100110011001100110011001100,
64'b1001100101100110100110010110011010011001011001101001100101100110,
64'b1100001111000011110000111100001100111100001111000011110000111100,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b0000111111110000000011111111000000001111111100000000111111110000,
64'b1111000000001111000011111111000011110000000011110000111111110000,
64'b1100001111000011110000111100001100111100001111000011110000111100,
64'b1111000000001111000011111111000011110000000011110000111111110000,
64'b1100110000110011110011000011001100110011110011000011001111001100,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b0011001100110011001100110011001111001100110011001100110011001100,
64'b0110011001100110100110011001100110011001100110010110011001100110,
64'b0011110011000011001111001100001111000011001111001100001100111100,
64'b1100110011001100001100110011001100110011001100111100110011001100,
64'b1100110011001100001100110011001100110011001100111100110011001100,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1111000011110000111100001111000011110000111100001111000011110000,
64'b0110100101101001011010010110100110010110100101101001011010010110,
64'b0101101010100101101001010101101001011010101001011010010101011010,
64'b1010010110100101101001011010010101011010010110100101101001011010,
64'b1010010110100101101001011010010101011010010110100101101001011010,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b0110011001100110100110011001100110011001100110010110011001100110,
64'b0101101001011010010110100101101001011010010110100101101001011010,
64'b1010101001010101010101011010101010101010010101010101010110101010,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b0101101010100101010110101010010110100101010110101010010101011010,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b0101101010100101101001010101101001011010101001011010010101011010,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1111111111111111000000000000000011111111111111110000000000000000,
64'b0101010110101010010101011010101001010101101010100101010110101010,
64'b0000111111110000111100000000111111110000000011110000111111110000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0011001111001100110011000011001111001100001100110011001111001100,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1111111111111111111111111111111100000000000000000000000000000000,
64'b0011001100110011110011001100110000110011001100111100110011001100,
64'b1111111100000000000000001111111100000000111111111111111100000000,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b0110100110010110011010011001011001101001100101100110100110010110,
64'b0011001111001100001100111100110000110011110011000011001111001100,
64'b0011001100110011001100110011001111001100110011001100110011001100,
64'b0011110011000011001111001100001111000011001111001100001100111100,
64'b1100001111000011001111000011110011000011110000110011110000111100,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b1010010110100101101001011010010101011010010110100101101001011010,
64'b1001011001101001011010011001011010010110011010010110100110010110,
64'b1100001111000011110000111100001100111100001111000011110000111100,
64'b1100001111000011001111000011110011000011110000110011110000111100,
64'b1001100101100110100110010110011010011001011001101001100101100110,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b1001100101100110100110010110011010011001011001101001100101100110,
64'b0110100110010110100101100110100110010110011010010110100110010110,
64'b0000111111110000000011111111000000001111111100000000111111110000,
64'b0101101010100101010110101010010110100101010110101010010101011010,
64'b1100001111000011001111000011110011000011110000110011110000111100,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b0101101010100101010110101010010110100101010110101010010101011010,
64'b0101101001011010101001011010010110100101101001010101101001011010,
64'b1001100101100110011001101001100101100110100110011001100101100110,
64'b0101010101010101101010101010101001010101010101011010101010101010,
64'b1001100101100110100110010110011010011001011001101001100101100110,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b0101010101010101010101010101010110101010101010101010101010101010,
64'b1111111111111111111111111111111100000000000000000000000000000000,
64'b1010010110100101010110100101101010100101101001010101101001011010,
64'b0000000011111111000000001111111111111111000000001111111100000000,
64'b0000000000000000111111111111111111111111111111110000000000000000,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b0101010110101010101010100101010110101010010101010101010110101010,
64'b0011001111001100001100111100110000110011110011000011001111001100,
64'b0101010110101010010101011010101001010101101010100101010110101010,
64'b0110011010011001100110010110011001100110100110011001100101100110,
64'b1001011010010110100101101001011010010110100101101001011010010110,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b1100110011001100001100110011001100110011001100111100110011001100,
64'b1010010110100101010110100101101010100101101001010101101001011010,
64'b0011001100110011110011001100110000110011001100111100110011001100,
64'b0011110000111100110000111100001111000011110000110011110000111100,
64'b1100001100111100110000110011110011000011001111001100001100111100,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000111100001111000011110000111111110000111100001111000011110000,
64'b0110011010011001011001101001100110011001011001101001100101100110,
64'b0000111100001111000011110000111111110000111100001111000011110000,
64'b1111000000001111111100000000111100001111111100000000111111110000,
64'b0101101010100101101001010101101001011010101001011010010101011010,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0101010110101010010101011010101001010101101010100101010110101010,
64'b0110100101101001100101101001011001101001011010011001011010010110,
64'b0101010110101010010101011010101001010101101010100101010110101010,
64'b1010101001010101010101011010101010101010010101010101010110101010,
64'b1001100101100110011001101001100101100110100110011001100101100110,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000011111111000000001111111111111111000000001111111100000000,
64'b1010010110100101101001011010010101011010010110100101101001011010,
64'b0000000000000000111111111111111111111111111111110000000000000000,
64'b0101010110101010101010100101010110101010010101010101010110101010,
64'b1111111111111111000000000000000011111111111111110000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0101010101010101101010101010101001010101010101011010101010101010,
64'b1001100101100110100110010110011010011001011001101001100101100110,
64'b0101010101010101010101010101010110101010101010101010101010101010,
64'b0110011001100110100110011001100110011001100110010110011001100110,
64'b0101010101010101010101010101010110101010101010101010101010101010,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0011001100110011001100110011001111001100110011001100110011001100,
64'b1100001111000011001111000011110011000011110000110011110000111100,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b0110100101101001011010010110100110010110100101101001011010010110,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b1111000011110000111100001111000011110000111100001111000011110000,
64'b0101101010100101010110101010010110100101010110101010010101011010,
64'b1111000011110000111100001111000011110000111100001111000011110000,
64'b1100001100111100110000110011110011000011001111001100001100111100,
64'b1001011010010110100101101001011010010110100101101001011010010110,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b1111111100000000111111110000000011111111000000001111111100000000,
64'b1100110000110011001100111100110011001100001100110011001111001100,
64'b0101010110101010010101011010101001010101101010100101010110101010,
64'b1111000000001111000011111111000011110000000011110000111111110000,
64'b1100001100111100110000110011110011000011001111001100001100111100,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1111111111111111000000000000000011111111111111110000000000000000,
64'b1111000011110000000011110000111100001111000011111111000011110000,
64'b0011001100110011110011001100110000110011001100111100110011001100,
64'b1111111100000000000000001111111100000000111111111111111100000000,
64'b1111000000001111000011111111000011110000000011110000111111110000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1100110000110011001100111100110011001100001100110011001111001100,
64'b1001100110011001100110011001100101100110011001100110011001100110,
64'b1001011010010110100101101001011010010110100101101001011010010110,
64'b1001100101100110011001101001100101100110100110011001100101100110,
64'b1001011001101001011010011001011010010110011010010110100110010110,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b1100001100111100110000110011110011000011001111001100001100111100,
64'b1010010101011010101001010101101010100101010110101010010101011010,
64'b0101101010100101010110101010010110100101010110101010010101011010,
64'b1010010101011010010110101010010101011010101001011010010101011010,
64'b1010101001010101010101011010101010101010010101010101010110101010,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b1111000000001111000011111111000011110000000011110000111111110000,
64'b1100110000110011001100111100110011001100001100110011001111001100,
64'b1100110000110011001100111100110011001100001100110011001111001100,
64'b1001100101100110011001101001100101100110100110011001100101100110,
64'b0110011001100110100110011001100110011001100110010110011001100110,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b1111111100000000000000001111111100000000111111111111111100000000,
64'b1111000011110000000011110000111100001111000011111111000011110000,
64'b1111000011110000000011110000111100001111000011111111000011110000,
64'b0011110000111100110000111100001111000011110000110011110000111100,
64'b0110100101101001011010010110100110010110100101101001011010010110,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b1001100101100110100110010110011010011001011001101001100101100110,
64'b0011001100110011001100110011001111001100110011001100110011001100,
64'b1001100101100110100110010110011010011001011001101001100101100110,
64'b1100001111000011110000111100001100111100001111000011110000111100,
64'b1010101001010101101010100101010101010101101010100101010110101010,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b0110100101101001100101101001011001101001011010011001011010010110,
64'b1111000011110000111100001111000011110000111100001111000011110000,
64'b0110100101101001100101101001011001101001011010011001011010010110,
64'b0000111111110000000011111111000000001111111100000000111111110000,
64'b1001100110011001011001100110011010011001100110010110011001100110,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b1001011001101001100101100110100101101001100101100110100110010110,
64'b1111111100000000111111110000000011111111000000001111111100000000,
64'b0011110011000011001111001100001111000011001111001100001100111100,
64'b0000000011111111111111110000000000000000111111111111111100000000,
64'b1100001111000011110000111100001100111100001111000011110000111100,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b1001011001101001011010011001011010010110011010010110100110010110,
64'b0101010101010101101010101010101001010101010101011010101010101010,
64'b1111000000001111000011111111000011110000000011110000111111110000,
64'b1010101010101010010101010101010101010101010101011010101010101010,
64'b0000111111110000000011111111000000001111111100000000111111110000,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b1100001100111100001111001100001100111100110000111100001100111100,
64'b0011001100110011001100110011001111001100110011001100110011001100,
64'b1111111100000000000000001111111100000000111111111111111100000000,
64'b0011001100110011001100110011001111001100110011001100110011001100,
64'b1010101001010101010101011010101010101010010101010101010110101010,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b1010010101011010010110101010010101011010101001011010010101011010,
64'b0101101001011010010110100101101001011010010110100101101001011010,
64'b1010101010101010010101010101010101010101010101011010101010101010,
64'b0101101001011010010110100101101001011010010110100101101001011010,
64'b0110011001100110100110011001100110011001100110010110011001100110,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000111100001111000011110000111111110000111100001111000011110000,
64'b1111000011110000000011110000111100001111000011111111000011110000,
64'b0011001100110011001100110011001111001100110011001100110011001100,
64'b0000111111110000111100000000111111110000000011110000111111110000,
64'b1111000000001111111100000000111100001111111100000000111111110000,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b0101101010100101010110101010010110100101010110101010010101011010,
64'b0101101010100101101001010101101001011010101001011010010101011010,
64'b0110100101101001011010010110100110010110100101101001011010010110,
64'b0101101001011010010110100101101001011010010110100101101001011010,
64'b0101101001011010101001011010010110100101101001010101101001011010,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b1100001100111100001111001100001100111100110000111100001100111100,
64'b0110100110010110011010011001011001101001100101100110100110010110,
64'b1111000000001111111100000000111100001111111100000000111111110000,
64'b1001011010010110011010010110100101101001011010011001011010010110,
64'b0011110000111100001111000011110000111100001111000011110000111100,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b1010010101011010010110101010010101011010101001011010010101011010,
64'b1001011001101001011010011001011010010110011010010110100110010110,
64'b0000000011111111111111110000000000000000111111111111111100000000,
64'b1001011001101001100101100110100101101001100101100110100110010110,
64'b1010010101011010101001010101101010100101010110101010010101011010,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b0011110011000011110000110011110000111100110000111100001100111100,
64'b1001100101100110100110010110011010011001011001101001100101100110,
64'b0011001100110011110011001100110000110011001100111100110011001100,
64'b0011001100110011001100110011001111001100110011001100110011001100,
64'b1001011010010110011010010110100101101001011010011001011010010110,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b0000000011111111111111110000000000000000111111111111111100000000,
64'b0011001100110011001100110011001111001100110011001100110011001100,
64'b0011110000111100001111000011110000111100001111000011110000111100,
64'b1111111100000000000000001111111100000000111111111111111100000000,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b0000000000000000111111111111111111111111111111110000000000000000,
64'b1111000011110000111100001111000011110000111100001111000011110000,
64'b1010010101011010101001010101101010100101010110101010010101011010,
64'b0000000000000000111111111111111111111111111111110000000000000000,
64'b1001011010010110100101101001011010010110100101101001011010010110,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b0101101001011010010110100101101001011010010110100101101001011010,
64'b1010010101011010010110101010010101011010101001011010010101011010,
64'b1111111100000000000000001111111100000000111111111111111100000000,
64'b1111000000001111000011111111000011110000000011110000111111110000,
64'b1001100110011001100110011001100101100110011001100110011001100110,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b0011110011000011001111001100001111000011001111001100001100111100,
64'b1100001100111100110000110011110011000011001111001100001100111100,
64'b1001100110011001011001100110011010011001100110010110011001100110,
64'b0101101001011010010110100101101001011010010110100101101001011010,
64'b1100110000110011110011000011001100110011110011000011001111001100,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b1111000000001111000011111111000011110000000011110000111111110000,
64'b0101101010100101101001010101101001011010101001011010010101011010,
64'b1100001111000011110000111100001100111100001111000011110000111100,
64'b0011001111001100001100111100110000110011110011000011001111001100,
64'b0000111100001111111100001111000000001111000011111111000011110000,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b0101101010100101101001010101101001011010101001011010010101011010,
64'b1100001100111100110000110011110011000011001111001100001100111100,
64'b0011110011000011001111001100001111000011001111001100001100111100,
64'b1010101001010101101010100101010101010101101010100101010110101010,
64'b1111000011110000111100001111000011110000111100001111000011110000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b1001011001101001011010011001011010010110011010010110100110010110,
64'b0000000011111111000000001111111111111111000000001111111100000000,
64'b1100001100111100001111001100001100111100110000111100001100111100,
64'b1001011001101001100101100110100101101001100101100110100110010110,
64'b1010010110100101101001011010010101011010010110100101101001011010,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b0110011010011001100110010110011001100110100110011001100101100110,
64'b0000111100001111000011110000111111110000111100001111000011110000,
64'b1001011001101001011010011001011010010110011010010110100110010110,
64'b1001100110011001100110011001100101100110011001100110011001100110,
64'b0110100101101001011010010110100110010110100101101001011010010110,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b0011110000111100110000111100001111000011110000110011110000111100,
64'b1111111100000000111111110000000011111111000000001111111100000000,
64'b0110100110010110100101100110100110010110011010010110100110010110,
64'b0011110000111100001111000011110000111100001111000011110000111100,
64'b0110100110010110011010011001011001101001100101100110100110010110,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b1111000000001111111100000000111100001111111100000000111111110000,
64'b0101010101010101101010101010101001010101010101011010101010101010,
64'b1100001100111100001111001100001100111100110000111100001100111100,
64'b1010010101011010101001010101101010100101010110101010010101011010,
64'b0011110011000011110000110011110000111100110000111100001100111100,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b1010101001010101010101011010101010101010010101010101010110101010,
64'b1001100110011001100110011001100101100110011001100110011001100110,
64'b0000111111110000111100000000111111110000000011110000111111110000,
64'b0110011010011001100110010110011001100110100110011001100101100110,
64'b0000111111110000111100000000111111110000000011110000111111110000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0110100101101001100101101001011001101001011010011001011010010110,
64'b1100110011001100001100110011001100110011001100111100110011001100,
64'b0110011010011001100110010110011001100110100110011001100101100110,
64'b1001100101100110100110010110011010011001011001101001100101100110,
64'b0000111100001111111100001111000000001111000011111111000011110000,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b1001011001101001100101100110100101101001100101100110100110010110,
64'b0000111100001111000011110000111111110000111100001111000011110000,
64'b1001011010010110011010010110100101101001011010011001011010010110,
64'b1100001111000011001111000011110011000011110000110011110000111100,
64'b0000000011111111000000001111111111111111000000001111111100000000,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b0011110011000011110000110011110000111100110000111100001100111100,
64'b0101010110101010010101011010101001010101101010100101010110101010,
64'b1001011001101001100101100110100101101001100101100110100110010110,
64'b0101101010100101010110101010010110100101010110101010010101011010,
64'b1111111111111111000000000000000011111111111111110000000000000000,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b1010010101011010010110101010010101011010101001011010010101011010,
64'b0011001100110011110011001100110000110011001100111100110011001100,
64'b0011110011000011110000110011110000111100110000111100001100111100,
64'b0110011010011001100110010110011001100110100110011001100101100110,
64'b0101010101010101010101010101010110101010101010101010101010101010,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b1001100101100110011001101001100101100110100110011001100101100110,
64'b1010010110100101101001011010010101011010010110100101101001011010,
64'b0000111111110000111100000000111111110000000011110000111111110000,
64'b0011110000111100110000111100001111000011110000110011110000111100,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b1001011010010110011010010110100101101001011010011001011010010110,
64'b1001100101100110100110010110011010011001011001101001100101100110,
64'b0101010110101010101010100101010110101010010101010101010110101010,
64'b0101101010100101010110101010010110100101010110101010010101011010,
64'b0101101001011010010110100101101001011010010110100101101001011010,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b1001100101100110100110010110011010011001011001101001100101100110,
64'b1001100110011001100110011001100101100110011001100110011001100110,
64'b1111111111111111000000000000000011111111111111110000000000000000,
64'b0110100101101001011010010110100110010110100101101001011010010110,
64'b0110100101101001011010010110100110010110100101101001011010010110,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b1100110011001100001100110011001100110011001100111100110011001100,
64'b1100110011001100001100110011001100110011001100111100110011001100,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b1100110011001100001100110011001100110011001100111100110011001100,
64'b1001100110011001100110011001100101100110011001100110011001100110,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b0000111100001111000011110000111111110000111100001111000011110000,
64'b1010010110100101101001011010010101011010010110100101101001011010,
64'b1001011010010110100101101001011010010110100101101001011010010110,
64'b0000111100001111000011110000111111110000111100001111000011110000,
64'b1001011010010110100101101001011010010110100101101001011010010110,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b1111111100000000111111110000000011111111000000001111111100000000,
64'b1001100101100110100110010110011010011001011001101001100101100110,
64'b0110100110010110011010011001011001101001100101100110100110010110,
64'b1111111100000000111111110000000011111111000000001111111100000000,
64'b0110100110010110011010011001011001101001100101100110100110010110,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b1111000011110000000011110000111100001111000011111111000011110000,
64'b0011001100110011001100110011001111001100110011001100110011001100,
64'b0000111111110000111100000000111111110000000011110000111111110000,
64'b1111000000001111111100000000111100001111111100000000111111110000,
64'b1100110011001100001100110011001100110011001100111100110011001100,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b1010101001010101101010100101010101010101101010100101010110101010,
64'b0101101001011010010110100101101001011010010110100101101001011010,
64'b0101010110101010101010100101010110101010010101010101010110101010,
64'b1010101001010101010101011010101010101010010101010101010110101010,
64'b1010010110100101101001011010010101011010010110100101101001011010,
64'b1010101010101010101010101010101010101010101010101010101010101010,
64'b0011001100110011110011001100110000110011001100111100110011001100,
64'b1001100101100110100110010110011010011001011001101001100101100110,
64'b1100110011001100001100110011001100110011001100111100110011001100,
64'b0110011001100110100110011001100110011001100110010110011001100110,
64'b0011001111001100001100111100110000110011110011000011001111001100,
64'b0110011001100110011001100110011001100110011001100110011001100110,
64'b0000111100001111000011110000111111110000111100001111000011110000,
64'b1100001111000011001111000011110011000011110000110011110000111100,
64'b0000111100001111000011110000111111110000111100001111000011110000,
64'b0110100101101001011010010110100110010110100101101001011010010110,
64'b1010010110100101010110100101101010100101101001010101101001011010,
64'b1100110011001100110011001100110011001100110011001100110011001100,
64'b0101010110101010010101011010101001010101101010100101010110101010,
64'b0101101010100101010110101010010110100101010110101010010101011010,
64'b1111111100000000111111110000000011111111000000001111111100000000,
64'b0110100110010110011010011001011001101001100101100110100110010110,
64'b0110011010011001011001101001100110011001011001101001100101100110,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0011001100110011110011001100110000110011001100111100110011001100,
64'b1100110000110011001100111100110011001100001100110011001111001100,
64'b0101010101010101101010101010101001010101010101011010101010101010,
64'b0011110011000011110000110011110000111100110000111100001100111100,
64'b1100001111000011001111000011110011000011110000110011110000111100,
64'b1010101010101010101010101010101010101010101010101010101010101010  


};
                                  
 

//*********************
//INNER SIGNAL DECLARATION
//*********************
//REGS
 wire [31:0]     crc_go_back_1    ;
wire         crc_en_go_back_1    ;
wire [MOD_WIDTH-1:0]      mod_go_back_1    ;

wire [31:0]     crc_go_back_2    ;
wire         crc_en_go_back_2    ;
wire [MOD_WIDTH-1:0]      mod_go_back_2    ;

wire [31:0]     crc_go_back_3    ;
wire         crc_en_go_back_3    ;
wire [MOD_WIDTH-1:0]      mod_go_back_3    ;

wire [31:0]     crc_go_back_4    ;
wire         crc_en_go_back_4    ;
wire [MOD_WIDTH-1:0]      mod_go_back_4    ;

wire [31:0]     crc_go_back_5    ;
wire         crc_en_go_back_5    ;
wire [MOD_WIDTH-1:0]      mod_go_back_5    ;

wire [31:0]     crc_go_back_6    ;
wire         crc_en_go_back_6    ;
wire [MOD_WIDTH-1:0]      mod_go_back_6    ;

wire [31:0]     crc_go_back_7    ;
wire         crc_en_go_back_7    ;
wire [MOD_WIDTH-1:0]      mod_go_back_7    ; 

//WIRES
 

//*********************
//INSTANTCE MODULE
//*********************


        go_back_stage    // 512
            # ( 
                    .MOD ( 7'd64 ) ,  // 128-64
                    .POLY ( POLY[6*32*64*6 +: 32*64*6] )  
                )
        go_back_stage_1  (     
            .clk             ( clk )   ,
            .rst             ( rst )   ,
            .crc             ( crc_in )   ,
            .crc_en          ( crc_en_in )   ,
            .mod             ( mod_in )   ,
            .crc_go_back     (    crc_go_back_1 )   ,
            .crc_en_go_back  ( crc_en_go_back_1 )   ,
            .mod_go_back     (    mod_go_back_1 )           
                      ) ;

        go_back_stage    // 256
            # ( 
                    .MOD ( 7'd32 ) , // 128-32
                    .POLY ( POLY[5*32*64*6 +: 32*64*6] )  
                )
        go_back_stage_2  (     
            .clk             ( clk )   ,
            .rst             ( rst )   ,
            .crc             ( crc_go_back_1 )   ,
            .crc_en          ( crc_en_go_back_1 )   ,
            .mod             ( mod_go_back_1 )   ,
            .crc_go_back     ( crc_go_back_2 )   ,
            .crc_en_go_back  ( crc_en_go_back_2 )   ,
            .mod_go_back     ( mod_go_back_2 )           
                      ) ;

        go_back_stage    // 128
            # ( 
                    .MOD ( 7'd16 ) , // 128-16
                    .POLY ( POLY[4*32*64*6 +: 32*64*6] )  
                )
        go_back_stage_3  (     
            .clk             ( clk )   ,
            .rst             ( rst )   ,
            .crc             ( crc_go_back_2 )   ,
            .crc_en          ( crc_en_go_back_2 )   ,
            .mod             ( mod_go_back_2 )   ,
            .crc_go_back     ( crc_go_back_3 )   ,
            .crc_en_go_back  ( crc_en_go_back_3 )   ,
            .mod_go_back     ( mod_go_back_3 )           
                      ) ;


        go_back_stage    // 64
            # ( 
                    .MOD ( 7'd8 ) , // 128-8
                    .POLY ( POLY[3*32*64*6 +: 32*64*6] )  
                )
        go_back_stage_4  (     
            .clk             ( clk )   ,
            .rst             ( rst )   ,
            .crc             ( crc_go_back_3 )   ,
            .crc_en          ( crc_en_go_back_3 )   ,
            .mod             ( mod_go_back_3 )   ,
            .crc_go_back     ( crc_go_back_4 )   ,
            .crc_en_go_back  ( crc_en_go_back_4 )   ,
            .mod_go_back     ( mod_go_back_4 )           
                      ) ;

        go_back_stage    // 32
            # ( 
                    .MOD ( 7'd4 ) , // 128-4
                    .POLY ( POLY[2*32*64*6 +: 32*64*6] )  
                )
        go_back_stage_5  (     
            .clk             ( clk )   ,
            .rst             ( rst )   ,
            .crc             ( crc_go_back_4 )   ,
            .crc_en          ( crc_en_go_back_4 )   ,
            .mod             ( mod_go_back_4 )   ,
            .crc_go_back     ( crc_go_back_5 )   ,
            .crc_en_go_back  ( crc_en_go_back_5 )   ,
            .mod_go_back     ( mod_go_back_5 )           
                      ) ;


        go_back_stage    // 16
            # ( 
                    .MOD ( 7'd2 ) , // 128-2
                    .POLY ( POLY[1*32*64*6 +: 32*64*6] )  
                )
        go_back_stage_6  (     
            .clk             ( clk )   ,
            .rst             ( rst )   ,
            .crc             ( crc_go_back_5 )   ,
            .crc_en          ( crc_en_go_back_5 )   ,
            .mod             ( mod_go_back_5 )   ,
            .crc_go_back     ( crc_go_back_6 )   ,
            .crc_en_go_back  ( crc_en_go_back_6 )   ,
            .mod_go_back     ( mod_go_back_6 )           
                      ) ;

        go_back_stage    // 8
            # ( 
                    .MOD ( 7'd1 ) , // 128-1
                    .POLY ( POLY[0 +: 32*64*6] )  
                )
        go_back_stage_7  (     
            .clk             ( clk )   ,
            .rst             ( rst )   ,
            .crc             ( crc_go_back_6 )   ,
            .crc_en          ( crc_en_go_back_6 )   ,
            .mod             ( mod_go_back_6 )   ,
            .crc_go_back     ( crc_out )   ,
            .crc_en_go_back  ( crc_out_en )   ,
            .mod_go_back     (  )           
                      ) ;


//*********************
//MAIN CORE
//********************* 





//*********************
endmodule   