
// **************************************************************
// COPYRIGHT(c)2015, Xidian University
// All rights reserved.
//
// IP LIB INDEX :  
// IP Name      :      
// File name    : 
// Module name  : 
// Full name    :  
//
// Author       : Liu-Huan 
// Email        : assasin9997@163.com 
// Data         : 
// Version      : V 1.0 
// 
// Abstract     : 
// Called by    :  
// 
// Modification history
// -----------------------------------------------------------------
// 
// 
//
// *****************************************************************

// *******************
// TIMESCALE
// ******************* 
`timescale 1ns/1ps 

// *******************
// INFORMATION
// *******************


//*******************
//DEFINE(s)
//*******************
//`define UDLY 1    //Unit delay, for non-blocking assignments in sequential logic


//*******************
//DEFINE MODULE PORT
//*******************
module  data_source_65   (     
            input 				clk     ,
            output  			sop     ,
            output  			eop     ,
            output  			dval    ,
            output  [2:0] 		mod     ,
            output  [63:0] 		dout         
              ) ;

//*******************
//DEFINE LOCAL PARAMETER
//*******************
//parameter(s)
                                    
 

//*********************
//INNER SIGNAL DECLARATION
//*********************
//REGS
  reg [79:0] mem [0:8191] ;
  reg [79:0] dout_ff = 80'b0 ;

//WIRES
 

//*********************
//INSTANTCE MODULE
//*********************

initial begin
mem[0]    = 80'h00000000000000000000;
mem[1]    = 80'h00000000000000000000;
mem[2]    = 80'h10100000010000010010;
mem[3]    = 80'h00109400000208004500;
mem[4]    = 80'h0010002f5efa0000fffd;
mem[5]    = 80'h0010da7ec0550102c000;
mem[6]    = 80'h00100001ffabffabffab;
mem[7]    = 80'h0010ff05c779b3610cfb;
mem[8]    = 80'h0010eb2114e13678f7a9;
mem[9]    = 80'h0010364f68afabc8ce69;
mem[10]   = 80'h01119000000000000000;
mem[11]   = 80'h10100000010000010010;
mem[12]   = 80'h00109400000208004500;
mem[13]   = 80'h0010002f5efb0000fffd;
mem[14]   = 80'h0010da7dc0550102c000;
mem[15]   = 80'h00100001ffabffabffab;
mem[16]   = 80'h0010ff04b6a79fb97539;
mem[17]   = 80'h001054eac666db8d27a9;
mem[18]   = 80'h0010673ea29a0ca699d0;
mem[19]   = 80'h01113600000000000000;
mem[20]   = 80'h00000000000000000000;
mem[21]   = 80'h00000000000000000000;
mem[22]   = 80'h00000000000000000000;
mem[23]   = 80'h10100000010000010010;
mem[24]   = 80'h00109400000208004500;
mem[25]   = 80'h0010002f5efc0000fffd;
mem[26]   = 80'h0010da7cc0550102c000;
mem[27]   = 80'h00100001ffabffabffab;
mem[28]   = 80'h0010ff039263756861b6;
mem[29]   = 80'h0010d4522977b7b1c6da;
mem[30]   = 80'h00108226f7fca0adbc2c;
mem[31]   = 80'h01118400000000000000;
mem[32]   = 80'h00000000000000000000;
mem[33]   = 80'h10100000010000010010;
mem[34]   = 80'h00109400000208004500;
mem[35]   = 80'h0010002f5efd0000fffd;
mem[36]   = 80'h0010da7bc0550102c000;
mem[37]   = 80'h00100001ffabffabffab;
mem[38]   = 80'h0010ff02e3bd59b01874;
mem[39]   = 80'h00106b99fbf05a44165b;
mem[40]   = 80'h0010d37f94716a42ac19;
mem[41]   = 80'h01116300000000000000;
mem[42]   = 80'h00000000000000000000;
mem[43]   = 80'h00000000000000000000;
mem[44]   = 80'h00000000000000000000;
mem[45]   = 80'h10100000010000010010;
mem[46]   = 80'h00109400000208004500;
mem[47]   = 80'h0010002f5efe0000fffd;
mem[48]   = 80'h0010da7ac0550102c000;
mem[49]   = 80'h00100001ffabffabffab;
mem[50]   = 80'h0010ff0171df2cd89233;
mem[51]   = 80'h0010abc58c786c5a66c8;
mem[52]   = 80'h001021b053024f541846;
mem[53]   = 80'h01112b00000000000000;
mem[54]   = 80'h00000000000000000000;
mem[55]   = 80'h00000000000000000000;
mem[56]   = 80'h00000000000000000000;
mem[57]   = 80'h10100000010000010010;
mem[58]   = 80'h00109400000208004500;
mem[59]   = 80'h0010002f5eff0000fffd;
mem[60]   = 80'h0010da79c0550102c000;
mem[61]   = 80'h00100001ffabffabffab;
mem[62]   = 80'h0010ff0000010000ebf1;
mem[63]   = 80'h0010140e5eff81afb6c9;
mem[64]   = 80'h001070f2a8934fd10b4d;
mem[65]   = 80'h01110300000000000000;
mem[66]   = 80'h00000000000000000000;
mem[67]   = 80'h10100000010000010010;
mem[68]   = 80'h00109400000208004500;
mem[69]   = 80'h0010002f5f000000fffd;
mem[70]   = 80'h0010da78c0550102c000;
mem[71]   = 80'h00100001ffabffabffab;
mem[72]   = 80'h0010ffff2f4b1bb73cb0;
mem[73]   = 80'h00108148ee82dafcf939;
mem[74]   = 80'h0010bf12303944980b45;
mem[75]   = 80'h01110200000000000000;
mem[76]   = 80'h00000000000000000000;
mem[77]   = 80'h00000000000000000000;
mem[78]   = 80'h00000000000000000000;
mem[79]   = 80'h10100000010000010010;
mem[80]   = 80'h00109400000208004500;
mem[81]   = 80'h0010002f5f010000fffd;
mem[82]   = 80'h0010da77c0550102c000;
mem[83]   = 80'h00100001ffabffabffab;
mem[84]   = 80'h0010fffe5e95376f4572;
mem[85]   = 80'h00103e833c05370928bb;
mem[86]   = 80'h0010ee2930142b3c7236;
mem[87]   = 80'h01116600000000000000;
mem[88]   = 80'h00000000000000000000;
mem[89]   = 80'h10100000010000010010;
mem[90]   = 80'h00109400000208004500;
mem[91]   = 80'h0010002f5f020000fffd;
mem[92]   = 80'h0010da76c0550102c000;
mem[93]   = 80'h00100001ffabffabffab;
mem[94]   = 80'h0010fffdccf74207cf35;
mem[95]   = 80'h0010fedf4b8d01175808;
mem[96]   = 80'h00101ce011614f52e640;
mem[97]   = 80'h0111f600000000000000;
mem[98]   = 80'h00000000000000000000;
mem[99]   = 80'h00000000000000000000;
mem[100]  = 80'h00000000000000000000;
mem[101]  = 80'h10100000010000010010;
mem[102]  = 80'h00109400000208004500;
mem[103]  = 80'h0010002f5f030000fffd;
mem[104]  = 80'h0010da75c0550102c000;
mem[105]  = 80'h00100001ffabffabffab;
mem[106]  = 80'h0010fffcbd296edfb6f7;
mem[107]  = 80'h00104114990aece28849;
mem[108]  = 80'h00104daf260859a6967d;
mem[109]  = 80'h01119300000000000000;
mem[110]  = 80'h00000000000000000000;
mem[111]  = 80'h10100000010000010010;
mem[112]  = 80'h00109400000208004500;
mem[113]  = 80'h0010002f5f040000fffd;
mem[114]  = 80'h0010da74c0550102c000;
mem[115]  = 80'h00100001ffabffabffab;
mem[116]  = 80'h0010fffb99ed840ea278;
mem[117]  = 80'h0010c1ac761b80de697a;
mem[118]  = 80'h0010a8babfb3b46cc44b;
mem[119]  = 80'h01117100000000000000;
mem[120]  = 80'h00000000000000000000;
mem[121]  = 80'h00000000000000000000;
mem[122]  = 80'h00000000000000000000;
mem[123]  = 80'h00000000000000000000;
mem[124]  = 80'h10100000010000010010;
mem[125]  = 80'h00109400000208004500;
mem[126]  = 80'h0010002f5f050000fffd;
mem[127]  = 80'h0010da73c0550102c000;
mem[128]  = 80'h00100001ffabffabffab;
mem[129]  = 80'h0010fffae833a8d6dbba;
mem[130]  = 80'h00107e67a49c6d2bb93b;
mem[131]  = 80'h0010f9f588dec64a8c95;
mem[132]  = 80'h01110200000000000000;
mem[133]  = 80'h10100000010000010010;
mem[134]  = 80'h00109400000208004500;
mem[135]  = 80'h0010002f5f060000fffd;
mem[136]  = 80'h0010da72c0550102c000;
mem[137]  = 80'h00100001ffabffabffab;
mem[138]  = 80'h0010fff97a51ddbe51fd;
mem[139]  = 80'h0010be3bd3145b35c968;
mem[140]  = 80'h00100b2c1bde783ec82a;
mem[141]  = 80'h01112600000000000000;
mem[142]  = 80'h00000000000000000000;
mem[143]  = 80'h00000000000000000000;
mem[144]  = 80'h00000000000000000000;
mem[145]  = 80'h10100000010000010010;
mem[146]  = 80'h00109400000208004500;
mem[147]  = 80'h0010002f5f070000fffd;
mem[148]  = 80'h0010da71c0550102c000;
mem[149]  = 80'h00100001ffabffabffab;
mem[150]  = 80'h0010fff80b8ff166283f;
mem[151]  = 80'h001001f00193b6c01928;
mem[152]  = 80'h00105a501d168fc1ec6d;
mem[153]  = 80'h01112f00000000000000;
mem[154]  = 80'h10100000010000010010;
mem[155]  = 80'h00109400000208004500;
mem[156]  = 80'h0010002f5f080000fffd;
mem[157]  = 80'h0010da70c0550102c000;
mem[158]  = 80'h00100001ffabffabffab;
mem[159]  = 80'h0010fff733d8081c78e2;
mem[160]  = 80'h0010bf4a0d36834c0b9e;
mem[161]  = 80'h0010c03cd2895c3c5d61;
mem[162]  = 80'h01111d00000000000000;
mem[163]  = 80'h00000000000000000000;
mem[164]  = 80'h00000000000000000000;
mem[165]  = 80'h00000000000000000000;
mem[166]  = 80'h10100000010000010010;
mem[167]  = 80'h00109400000208004500;
mem[168]  = 80'h0010002f5f090000fffd;
mem[169]  = 80'h0010da6fc0550102c000;
mem[170]  = 80'h00100001ffabffabffab;
mem[171]  = 80'h0010fff6420624c40120;
mem[172]  = 80'h00100081dfb16eb9dbdf;
mem[173]  = 80'h00109173e5def54d13f6;
mem[174]  = 80'h0111cb00000000000000;
mem[175]  = 80'h00000000000000000000;
mem[176]  = 80'h10100000010000010010;
mem[177]  = 80'h00109400000208004500;
mem[178]  = 80'h0010002f5f0a0000fffd;
mem[179]  = 80'h0010da6ec0550102c000;
mem[180]  = 80'h00100001ffabffabffab;
mem[181]  = 80'h0010fff5d06451ac8b67;
mem[182]  = 80'h0010c0dda83958a7ab6c;
mem[183]  = 80'h001063bac4abbc56db5f;
mem[184]  = 80'h01111e00000000000000;
mem[185]  = 80'h00000000000000000000;
mem[186]  = 80'h00000000000000000000;
mem[187]  = 80'h00000000000000000000;
mem[188]  = 80'h00000000000000000000;
mem[189]  = 80'h10100000010000010010;
mem[190]  = 80'h00109400000208004500;
mem[191]  = 80'h0010002f5f0b0000fffd;
mem[192]  = 80'h0010da6dc0550102c000;
mem[193]  = 80'h00100001ffabffabffab;
mem[194]  = 80'h0010fff4a1ba7d74f2a5;
mem[195]  = 80'h00107f167abeb55274ed;
mem[196]  = 80'h001032cf9652001d140a;
mem[197]  = 80'h01110a00000000000000;
mem[198]  = 80'h00000000000000000000;
mem[199]  = 80'h10100000010000010010;
mem[200]  = 80'h00109400000208004500;
mem[201]  = 80'h0010002f5f0c0000fffd;
mem[202]  = 80'h0010da6cc0550102c000;
mem[203]  = 80'h00100001ffabffabffab;
mem[204]  = 80'h0010fff3857e97a5e62a;
mem[205]  = 80'h0010ffae95afd96e959e;
mem[206]  = 80'h0010d7d7c3795c42f29c;
mem[207]  = 80'h01114000000000000000;
mem[208]  = 80'h00000000000000000000;
mem[209]  = 80'h00000000000000000000;
mem[210]  = 80'h00000000000000000000;
mem[211]  = 80'h10100000010000010010;
mem[212]  = 80'h00109400000208004500;
mem[213]  = 80'h0010002f5f0d0000fffd;
mem[214]  = 80'h0010da6bc0550102c000;
mem[215]  = 80'h00100001ffabffabffab;
mem[216]  = 80'h0010fff2f4a0bb7d9fe8;
mem[217]  = 80'h001040654728349b4598;
mem[218]  = 80'h0010860caf38787da8ed;
mem[219]  = 80'h0111c800000000000000;
mem[220]  = 80'h00000000000000000000;
mem[221]  = 80'h10100000010000010010;
mem[222]  = 80'h00109400000208004500;
mem[223]  = 80'h0010002f5f0e0000fffd;
mem[224]  = 80'h0010da6ac0550102c000;
mem[225]  = 80'h00100001ffabffabffab;
mem[226]  = 80'h0010fff166c2ce1515af;
mem[227]  = 80'h0010803930a002853513;
mem[228]  = 80'h00107449b2cba5419828;
mem[229]  = 80'h0111e500000000000000;
mem[230]  = 80'h00000000000000000000;
mem[231]  = 80'h10100000010000010010;
mem[232]  = 80'h00109400000208004500;
mem[233]  = 80'h0010002f5f0f0000fffd;
mem[234]  = 80'h0010da69c0550102c000;
mem[235]  = 80'h00100001ffabffabffab;
mem[236]  = 80'h0010fff0171ce2cd6c6d;
mem[237]  = 80'h00103ff2e227ef70e58a;
mem[238]  = 80'h0010259a0b08719ee9c7;
mem[239]  = 80'h01114300000000000000;
mem[240]  = 80'h00000000000000000000;
mem[241]  = 80'h00000000000000000000;
mem[242]  = 80'h00000000000000000000;
mem[243]  = 80'h10100000010000010010;
mem[244]  = 80'h00109400000208004500;
mem[245]  = 80'h0010002f5f100000fffd;
mem[246]  = 80'h0010da68c0550102c000;
mem[247]  = 80'h00100001ffabffabffab;
mem[248]  = 80'h0010ffef166d3ce1b414;
mem[249]  = 80'h0010fd4d29ea699d107e;
mem[250]  = 80'h001040902cc9e9602356;
mem[251]  = 80'h0111d400000000000000;
mem[252]  = 80'h00000000000000000000;
mem[253]  = 80'h10100000010000010010;
mem[254]  = 80'h00109400000208004500;
mem[255]  = 80'h0010002f5f110000fffd;
mem[256]  = 80'h0010da67c0550102c000;
mem[257]  = 80'h00100001ffabffabffab;
mem[258]  = 80'h0010ffee67b31039cdd6;
mem[259]  = 80'h00104286fb6d8468c077;
mem[260]  = 80'h0010115b7e1ea77b4041;
mem[261]  = 80'h01112900000000000000;
mem[262]  = 80'h00000000000000000000;
mem[263]  = 80'h00000000000000000000;
mem[264]  = 80'h00000000000000000000;
mem[265]  = 80'h10100000010000010010;
mem[266]  = 80'h00109400000208004500;
mem[267]  = 80'h0010002f5f120000fffd;
mem[268]  = 80'h0010da66c0550102c000;
mem[269]  = 80'h00100001ffabffabffab;
mem[270]  = 80'h0010ffedf5d165514791;
mem[271]  = 80'h001082da8ce5b276b0fc;
mem[272]  = 80'h0010e31e630ba35d4eaf;
mem[273]  = 80'h0111f300000000000000;
mem[274]  = 80'h00000000000000000000;
mem[275]  = 80'h10100000010000010010;
mem[276]  = 80'h00109400000208004500;
mem[277]  = 80'h0010002f5f130000fffd;
mem[278]  = 80'h0010da65c0550102c000;
mem[279]  = 80'h00100001ffabffabffab;
mem[280]  = 80'h0010ffec840f49893e53;
mem[281]  = 80'h00103d115e625f836085;
mem[282]  = 80'h0010b2dd68cd7c2c7462;
mem[283]  = 80'h01113f00000000000000;
mem[284]  = 80'h00000000000000000000;
mem[285]  = 80'h00000000000000000000;
mem[286]  = 80'h00000000000000000000;
mem[287]  = 80'h00000000000000000000;
mem[288]  = 80'h10100000010000010010;
mem[289]  = 80'h00109400000208004500;
mem[290]  = 80'h0010002f5f140000fffd;
mem[291]  = 80'h0010da64c0550102c000;
mem[292]  = 80'h00100001ffabffabffab;
mem[293]  = 80'h0010ffeba0cba3582adc;
mem[294]  = 80'h0010bda9b17333bf803f;
mem[295]  = 80'h0010575ec19954b6ea34;
mem[296]  = 80'h0111cc00000000000000;
mem[297]  = 80'h10100000010000010010;
mem[298]  = 80'h00109400000208004500;
mem[299]  = 80'h0010002f5f150000fffd;
mem[300]  = 80'h0010da63c0550102c000;
mem[301]  = 80'h00100001ffabffabffab;
mem[302]  = 80'h0010ffead1158f80531e;
mem[303]  = 80'h0010026263f4de4a5076;
mem[304]  = 80'h001006985fb150ead029;
mem[305]  = 80'h01112100000000000000;
mem[306]  = 80'h00000000000000000000;
mem[307]  = 80'h00000000000000000000;
mem[308]  = 80'h00000000000000000000;
mem[309]  = 80'h10100000010000010010;
mem[310]  = 80'h00109400000208004500;
mem[311]  = 80'h0010002f5f160000fffd;
mem[312]  = 80'h0010da62c0550102c000;
mem[313]  = 80'h00100001ffabffabffab;
mem[314]  = 80'h0010ffe94377fae8d959;
mem[315]  = 80'h0010c23e147ce85420bd;
mem[316]  = 80'h0010f4d08ebe84564bbe;
mem[317]  = 80'h0111a800000000000000;
mem[318]  = 80'h00000000000000000000;
mem[319]  = 80'h10100000010000010010;
mem[320]  = 80'h00109400000208004500;
mem[321]  = 80'h0010002f5f170000fffd;
mem[322]  = 80'h0010da61c0550102c000;
mem[323]  = 80'h00100001ffabffabffab;
mem[324]  = 80'h0010ffe832a9d630a09b;
mem[325]  = 80'h00107df5c6fb05a1f0e4;
mem[326]  = 80'h0010a515631512016b88;
mem[327]  = 80'h01113400000000000000;
mem[328]  = 80'h00000000000000000000;
mem[329]  = 80'h00000000000000000000;
mem[330]  = 80'h00000000000000000000;
mem[331]  = 80'h10100000010000010010;
mem[332]  = 80'h00109400000208004500;
mem[333]  = 80'h0010002f5f180000fffd;
mem[334]  = 80'h0010da60c0550102c000;
mem[335]  = 80'h00100001ffabffabffab;
mem[336]  = 80'h0010ffe70afe2f4af046;
mem[337]  = 80'h0010c34fca5e302de2da;
mem[338]  = 80'h00103feb9de756ccf9bf;
mem[339]  = 80'h01117800000000000000;
mem[340]  = 80'h00000000000000000000;
mem[341]  = 80'h10100000010000010010;
mem[342]  = 80'h00109400000208004500;
mem[343]  = 80'h0010002f5f190000fffd;
mem[344]  = 80'h0010da5fc0550102c000;
mem[345]  = 80'h00100001ffabffabffab;
mem[346]  = 80'h0010ffe67b2003928984;
mem[347]  = 80'h00107c8418d9ddd83293;
mem[348]  = 80'h00106e2d03ebdf20cc51;
mem[349]  = 80'h01117f00000000000000;
mem[350]  = 80'h00000000000000000000;
mem[351]  = 80'h00000000000000000000;
mem[352]  = 80'h00000000000000000000;
mem[353]  = 80'h00000000000000000000;
mem[354]  = 80'h10100000010000010010;
mem[355]  = 80'h00109400000208004500;
mem[356]  = 80'h0010002f5f1a0000fffd;
mem[357]  = 80'h0010da5ec0550102c000;
mem[358]  = 80'h00100001ffabffabffab;
mem[359]  = 80'h0010ffe5e94276fa03c3;
mem[360]  = 80'h0010bcd86f51ebc6425b;
mem[361]  = 80'h00109c30819d230e2033;
mem[362]  = 80'h01112900000000000000;
mem[363]  = 80'h10100000010000010010;
mem[364]  = 80'h00109400000208004500;
mem[365]  = 80'h0010002f5f1b0000fffd;
mem[366]  = 80'h0010da5dc0550102c000;
mem[367]  = 80'h00100001ffabffabffab;
mem[368]  = 80'h0010ffe4989c5a227a01;
mem[369]  = 80'h00100313bdd606339222;
mem[370]  = 80'h0010cdf38a27e15c4072;
mem[371]  = 80'h01110500000000000000;
mem[372]  = 80'h00000000000000000000;
mem[373]  = 80'h00000000000000000000;
mem[374]  = 80'h00000000000000000000;
mem[375]  = 80'h10100000010000010010;
mem[376]  = 80'h00109400000208004500;
mem[377]  = 80'h0010002f5f1c0000fffd;
mem[378]  = 80'h0010da5cc0550102c000;
mem[379]  = 80'h00100001ffabffabffab;
mem[380]  = 80'h0010ffe3bc58b0f36e8e;
mem[381]  = 80'h001083ab52c76a0f7359;
mem[382]  = 80'h001028627603d18c8ad3;
mem[383]  = 80'h01112600000000000000;
mem[384]  = 80'h00000000000000000000;
mem[385]  = 80'h10100000010000010010;
mem[386]  = 80'h00109400000208004500;
mem[387]  = 80'h0010002f5f1d0000fffd;
mem[388]  = 80'h0010da5bc0550102c000;
mem[389]  = 80'h00100001ffabffabffab;
mem[390]  = 80'h0010ffe2cd869c2b174c;
mem[391]  = 80'h00103c60804087faa0d0;
mem[392]  = 80'h001079ebecc732759f15;
mem[393]  = 80'h0111e300000000000000;
mem[394]  = 80'h00000000000000000000;
mem[395]  = 80'h00000000000000000000;
mem[396]  = 80'h00000000000000000000;
mem[397]  = 80'h10100000010000010010;
mem[398]  = 80'h00109400000208004500;
mem[399]  = 80'h0010002f5f1e0000fffd;
mem[400]  = 80'h0010da5ac0550102c000;
mem[401]  = 80'h00100001ffabffabffab;
mem[402]  = 80'h0010ffe15fe4e9439d0b;
mem[403]  = 80'h0010fc3cf7c8b1e4d05b;
mem[404]  = 80'h00108baef1f525e86280;
mem[405]  = 80'h01116700000000000000;
mem[406]  = 80'h00000000000000000000;
mem[407]  = 80'h00000000000000000000;
mem[408]  = 80'h00000000000000000000;
mem[409]  = 80'h10100000010000010010;
mem[410]  = 80'h00109400000208004500;
mem[411]  = 80'h0010002f5f1f0000fffd;
mem[412]  = 80'h0010da59c0550102c000;
mem[413]  = 80'h00100001ffabffabffab;
mem[414]  = 80'h0010ffe02e3ac59be4c9;
mem[415]  = 80'h001043f7254f5c110042;
mem[416]  = 80'h0010da66d07eb6072fdf;
mem[417]  = 80'h01117b00000000000000;
mem[418]  = 80'h00000000000000000000;
mem[419]  = 80'h10100000010000010010;
mem[420]  = 80'h00109400000208004500;
mem[421]  = 80'h0010002f5f200000fffd;
mem[422]  = 80'h0010da58c0550102c000;
mem[423]  = 80'h00100001ffabffabffab;
mem[424]  = 80'h0010ffdf5d07551a2df8;
mem[425]  = 80'h001079436053bc3f3ba2;
mem[426]  = 80'h0010418afd030f0a61a3;
mem[427]  = 80'h0111dd00000000000000;
mem[428]  = 80'h00000000000000000000;
mem[429]  = 80'h00000000000000000000;
mem[430]  = 80'h00000000000000000000;
mem[431]  = 80'h10100000010000010010;
mem[432]  = 80'h00109400000208004500;
mem[433]  = 80'h0010002f5f210000fffd;
mem[434]  = 80'h0010da57c0550102c000;
mem[435]  = 80'h00100001ffabffabffab;
mem[436]  = 80'h0010ffde2cd979c2543a;
mem[437]  = 80'h0010c688b2d451caeb2b;
mem[438]  = 80'h0010105a379e06a35c32;
mem[439]  = 80'h0111a800000000000000;
mem[440]  = 80'h00000000000000000000;
mem[441]  = 80'h10100000010000010010;
mem[442]  = 80'h00109400000208004500;
mem[443]  = 80'h0010002f5f220000fffd;
mem[444]  = 80'h0010da56c0550102c000;
mem[445]  = 80'h00100001ffabffabffab;
mem[446]  = 80'h0010ffddbebb0caade7d;
mem[447]  = 80'h001006d4c55c67d49ba0;
mem[448]  = 80'h0010e21f2a79790e7981;
mem[449]  = 80'h01119300000000000000;
mem[450]  = 80'h00000000000000000000;
mem[451]  = 80'h00000000000000000000;
mem[452]  = 80'h00000000000000000000;
mem[453]  = 80'h10100000010000010010;
mem[454]  = 80'h00109400000208004500;
mem[455]  = 80'h0010002f5f230000fffd;
mem[456]  = 80'h0010da55c0550102c000;
mem[457]  = 80'h00100001ffabffabffab;
mem[458]  = 80'h0010ffdccf652072a7bf;
mem[459]  = 80'h0010b91f17db8a214bd9;
mem[460]  = 80'h0010b3dc21b9ebd4d97b;
mem[461]  = 80'h01110100000000000000;
mem[462]  = 80'h00000000000000000000;
mem[463]  = 80'h10100000010000010010;
mem[464]  = 80'h00109400000208004500;
mem[465]  = 80'h0010002f5f240000fffd;
mem[466]  = 80'h0010da54c0550102c000;
mem[467]  = 80'h00100001ffabffabffab;
mem[468]  = 80'h0010ffdbeba1caa3b330;
mem[469]  = 80'h001039a7f8cae61daae2;
mem[470]  = 80'h0010564011fb6aaae19c;
mem[471]  = 80'h0111c800000000000000;
mem[472]  = 80'h00000000000000000000;
mem[473]  = 80'h00000000000000000000;
mem[474]  = 80'h00000000000000000000;
mem[475]  = 80'h00000000000000000000;
mem[476]  = 80'h10100000010000010010;
mem[477]  = 80'h00109400000208004500;
mem[478]  = 80'h0010002f5f250000fffd;
mem[479]  = 80'h0010da53c0550102c000;
mem[480]  = 80'h00100001ffabffabffab;
mem[481]  = 80'h0010ffda9a7fe67bcaf2;
mem[482]  = 80'h0010866c2a4d0be87aab;
mem[483]  = 80'h001007868f63e5e62f2e;
mem[484]  = 80'h0111bb00000000000000;
mem[485]  = 80'h10100000010000010010;
mem[486]  = 80'h00109400000208004500;
mem[487]  = 80'h0010002f5f260000fffd;
mem[488]  = 80'h0010da52c0550102c000;
mem[489]  = 80'h00100001ffabffabffab;
mem[490]  = 80'h0010ffd9081d931340b5;
mem[491]  = 80'h001046305dc53df60be7;
mem[492]  = 80'h0010f57b61f1de358cba;
mem[493]  = 80'h01116600000000000000;
mem[494]  = 80'h00000000000000000000;
mem[495]  = 80'h00000000000000000000;
mem[496]  = 80'h00000000000000000000;
mem[497]  = 80'h10100000010000010010;
mem[498]  = 80'h00109400000208004500;
mem[499]  = 80'h0010002f5f270000fffd;
mem[500]  = 80'h0010da51c0550102c000;
mem[501]  = 80'h00100001ffabffabffab;
mem[502]  = 80'h0010ffd879c3bfcb3977;
mem[503]  = 80'h0010f9fb8f42d003dba6;
mem[504]  = 80'h0010a43456035ddbc857;
mem[505]  = 80'h01111100000000000000;
mem[506]  = 80'h10100000010000010010;
mem[507]  = 80'h00109400000208004500;
mem[508]  = 80'h0010002f5f280000fffd;
mem[509]  = 80'h0010da50c0550102c000;
mem[510]  = 80'h00100001ffabffabffab;
mem[511]  = 80'h0010ffd7419446b169aa;
mem[512]  = 80'h0010474183e7e58fc900;
mem[513]  = 80'h00103e5bea236bdaa6b2;
mem[514]  = 80'h0111d700000000000000;
mem[515]  = 80'h00000000000000000000;
mem[516]  = 80'h00000000000000000000;
mem[517]  = 80'h00000000000000000000;
mem[518]  = 80'h10100000010000010010;
mem[519]  = 80'h00109400000208004500;
mem[520]  = 80'h0010002f5f290000fffd;
mem[521]  = 80'h0010da4fc0550102c000;
mem[522]  = 80'h00100001ffabffabffab;
mem[523]  = 80'h0010ffd6304a6a691068;
mem[524]  = 80'h0010f88a5160087a1941;
mem[525]  = 80'h00106f14dd529c7c1728;
mem[526]  = 80'h01114e00000000000000;
mem[527]  = 80'h00000000000000000000;
mem[528]  = 80'h10100000010000010010;
mem[529]  = 80'h00109400000208004500;
mem[530]  = 80'h0010002f5f2a0000fffd;
mem[531]  = 80'h0010da4ec0550102c000;
mem[532]  = 80'h00100001ffabffabffab;
mem[533]  = 80'h0010ffd5a2281f019a2f;
mem[534]  = 80'h001038d626e83e646902;
mem[535]  = 80'h00109dce3dddc1321f5b;
mem[536]  = 80'h0111a800000000000000;
mem[537]  = 80'h00000000000000000000;
mem[538]  = 80'h00000000000000000000;
mem[539]  = 80'h00000000000000000000;
mem[540]  = 80'h00000000000000000000;
mem[541]  = 80'h10100000010000010010;
mem[542]  = 80'h00109400000208004500;
mem[543]  = 80'h0010002f5f2b0000fffd;
mem[544]  = 80'h0010da4dc0550102c000;
mem[545]  = 80'h00100001ffabffabffab;
mem[546]  = 80'h0010ffd4d3f633d9e3ed;
mem[547]  = 80'h0010871df46fd391b943;
mem[548]  = 80'h0010cc810a8934ba948d;
mem[549]  = 80'h01119e00000000000000;
mem[550]  = 80'h00000000000000000000;
mem[551]  = 80'h10100000010000010010;
mem[552]  = 80'h00109400000208004500;
mem[553]  = 80'h0010002f5f2c0000fffd;
mem[554]  = 80'h0010da4cc0550102c000;
mem[555]  = 80'h00100001ffabffabffab;
mem[556]  = 80'h0010ffd3f732d908f762;
mem[557]  = 80'h001007a51b7ebfad5800;
mem[558]  = 80'h0010299cca2009665467;
mem[559]  = 80'h01112f00000000000000;
mem[560]  = 80'h00000000000000000000;
mem[561]  = 80'h00000000000000000000;
mem[562]  = 80'h00000000000000000000;
mem[563]  = 80'h10100000010000010010;
mem[564]  = 80'h00109400000208004500;
mem[565]  = 80'h0010002f5f2d0000fffd;
mem[566]  = 80'h0010da4bc0550102c000;
mem[567]  = 80'h00100001ffabffabffab;
mem[568]  = 80'h0010ffd286ecf5d08ea0;
mem[569]  = 80'h0010b86ec9f952588800;
mem[570]  = 80'h001078ed00211ee41bc5;
mem[571]  = 80'h0111c100000000000000;
mem[572]  = 80'h00000000000000000000;
mem[573]  = 80'h10100000010000010010;
mem[574]  = 80'h00109400000208004500;
mem[575]  = 80'h0010002f5f2e0000fffd;
mem[576]  = 80'h0010da4ac0550102c000;
mem[577]  = 80'h00100001ffabffabffab;
mem[578]  = 80'h0010ffd1148e80b804e7;
mem[579]  = 80'h00107832be716446f883;
mem[580]  = 80'h00108a21b4709374b9f1;
mem[581]  = 80'h0111b100000000000000;
mem[582]  = 80'h00000000000000000000;
mem[583]  = 80'h10100000010000010010;
mem[584]  = 80'h00109400000208004500;
mem[585]  = 80'h0010002f5f2f0000fffd;
mem[586]  = 80'h0010da49c0550102c000;
mem[587]  = 80'h00100001ffabffabffab;
mem[588]  = 80'h0010ffd06550ac607d25;
mem[589]  = 80'h0010c7f96cf689b32f02;
mem[590]  = 80'h0010dbfd47b55f435164;
mem[591]  = 80'h01115d00000000000000;
mem[592]  = 80'h00000000000000000000;
mem[593]  = 80'h00000000000000000000;
mem[594]  = 80'h00000000000000000000;
mem[595]  = 80'h10100000010000010010;
mem[596]  = 80'h00109400000208004500;
mem[597]  = 80'h0010002f5f300000fffd;
mem[598]  = 80'h0010da48c0550102c000;
mem[599]  = 80'h00100001ffabffabffab;
mem[600]  = 80'h0010ffcf6421724ca55c;
mem[601]  = 80'h00100546a73b0f5edaee;
mem[602]  = 80'h0010be7dba19742e0ab1;
mem[603]  = 80'h0111a500000000000000;
mem[604]  = 80'h00000000000000000000;
mem[605]  = 80'h10100000010000010010;
mem[606]  = 80'h00109400000208004500;
mem[607]  = 80'h0010002f5f310000fffd;
mem[608]  = 80'h0010da47c0550102c000;
mem[609]  = 80'h00100001ffabffabffab;
mem[610]  = 80'h0010ffce15ff5e94dc9e;
mem[611]  = 80'h0010ba8d75bce2ab0aef;
mem[612]  = 80'h0010ef3f41da5f84367b;
mem[613]  = 80'h0111e100000000000000;
mem[614]  = 80'h00000000000000000000;
mem[615]  = 80'h00000000000000000000;
mem[616]  = 80'h00000000000000000000;
mem[617]  = 80'h10100000010000010010;
mem[618]  = 80'h00109400000208004500;
mem[619]  = 80'h0010002f5f320000fffd;
mem[620]  = 80'h0010da46c0550102c000;
mem[621]  = 80'h00100001ffabffabffab;
mem[622]  = 80'h0010ffcd879d2bfc56d9;
mem[623]  = 80'h00107ad10234d4b57a6c;
mem[624]  = 80'h00101df3f5a4156afb53;
mem[625]  = 80'h01118600000000000000;
mem[626]  = 80'h00000000000000000000;
mem[627]  = 80'h10100000010000010010;
mem[628]  = 80'h00109400000208004500;
mem[629]  = 80'h0010002f5f330000fffd;
mem[630]  = 80'h0010da45c0550102c000;
mem[631]  = 80'h00100001ffabffabffab;
mem[632]  = 80'h0010ffccf64307242f1b;
mem[633]  = 80'h0010c51ad0b33940aaee;
mem[634]  = 80'h00104cffc5b346b5e7f6;
mem[635]  = 80'h01114f00000000000000;
mem[636]  = 80'h00000000000000000000;
mem[637]  = 80'h00000000000000000000;
mem[638]  = 80'h00000000000000000000;
mem[639]  = 80'h00000000000000000000;
mem[640]  = 80'h10100000010000010010;
mem[641]  = 80'h00109400000208004500;
mem[642]  = 80'h0010002f5f340000fffd;
mem[643]  = 80'h0010da44c0550102c000;
mem[644]  = 80'h00100001ffabffabffab;
mem[645]  = 80'h0010ffcbd287edf53b94;
mem[646]  = 80'h001045a23fa2557c4bad;
mem[647]  = 80'h0010a9e205d22dee8e37;
mem[648]  = 80'h01117f00000000000000;
mem[649]  = 80'h10100000010000010010;
mem[650]  = 80'h00109400000208004500;
mem[651]  = 80'h0010002f5f350000fffd;
mem[652]  = 80'h0010da43c0550102c000;
mem[653]  = 80'h00100001ffabffabffab;
mem[654]  = 80'h0010ffcaa359c12d4256;
mem[655]  = 80'h0010fa69ed25b8899bec;
mem[656]  = 80'h0010f8ad32a3f17a15f0;
mem[657]  = 80'h0111db00000000000000;
mem[658]  = 80'h00000000000000000000;
mem[659]  = 80'h00000000000000000000;
mem[660]  = 80'h00000000000000000000;
mem[661]  = 80'h10100000010000010010;
mem[662]  = 80'h00109400000208004500;
mem[663]  = 80'h0010002f5f360000fffd;
mem[664]  = 80'h0010da42c0550102c000;
mem[665]  = 80'h00100001ffabffabffab;
mem[666]  = 80'h0010ffc9313bb445c811;
mem[667]  = 80'h00103a359aad8e97eb2f;
mem[668]  = 80'h00100a6c4a8daebedc39;
mem[669]  = 80'h01110e00000000000000;
mem[670]  = 80'h00000000000000000000;
mem[671]  = 80'h10100000010000010010;
mem[672]  = 80'h00109400000208004500;
mem[673]  = 80'h0010002f5f370000fffd;
mem[674]  = 80'h0010da41c0550102c000;
mem[675]  = 80'h00100001ffabffabffab;
mem[676]  = 80'h0010ffc840e5989db1d3;
mem[677]  = 80'h001085fe482a63623b6e;
mem[678]  = 80'h00105b237dc42e99beec;
mem[679]  = 80'h0111e700000000000000;
mem[680]  = 80'h00000000000000000000;
mem[681]  = 80'h00000000000000000000;
mem[682]  = 80'h00000000000000000000;
mem[683]  = 80'h10100000010000010010;
mem[684]  = 80'h00109400000208004500;
mem[685]  = 80'h0010002f5f380000fffd;
mem[686]  = 80'h0010da40c0550102c000;
mem[687]  = 80'h00100001ffabffabffab;
mem[688]  = 80'h0010ffc778b261e7e10e;
mem[689]  = 80'h00103b44448f56ee2848;
mem[690]  = 80'h0010c16069251a8954ae;
mem[691]  = 80'h01119800000000000000;
mem[692]  = 80'h00000000000000000000;
mem[693]  = 80'h10100000010000010010;
mem[694]  = 80'h00109400000208004500;
mem[695]  = 80'h0010002f5f390000fffd;
mem[696]  = 80'h0010da3fc0550102c000;
mem[697]  = 80'h00100001ffabffabffab;
mem[698]  = 80'h0010ffc6096c4d3f98cc;
mem[699]  = 80'h0010848f9608bb1bf808;
mem[700]  = 80'h0010901c6fe842a4f652;
mem[701]  = 80'h01112900000000000000;
mem[702]  = 80'h00000000000000000000;
mem[703]  = 80'h00000000000000000000;
mem[704]  = 80'h00000000000000000000;
mem[705]  = 80'h00000000000000000000;
mem[706]  = 80'h10100000010000010010;
mem[707]  = 80'h00109400000208004500;
mem[708]  = 80'h0010002f5f3a0000fffd;
mem[709]  = 80'h0010da3ec0550102c000;
mem[710]  = 80'h00100001ffabffabffab;
mem[711]  = 80'h0010ffc59b0e3857128b;
mem[712]  = 80'h001044d3e1808d0588cb;
mem[713]  = 80'h001062dd17476351cabe;
mem[714]  = 80'h01116900000000000000;
mem[715]  = 80'h10100000010000010010;
mem[716]  = 80'h00109400000208004500;
mem[717]  = 80'h0010002f5f3b0000fffd;
mem[718]  = 80'h0010da3dc0550102c000;
mem[719]  = 80'h00100001ffabffabffab;
mem[720]  = 80'h0010ffc4ead0148f6b49;
mem[721]  = 80'h0010fb18330760f0588a;
mem[722]  = 80'h001033922065598840d6;
mem[723]  = 80'h01112d00000000000000;
mem[724]  = 80'h00000000000000000000;
mem[725]  = 80'h00000000000000000000;
mem[726]  = 80'h00000000000000000000;
mem[727]  = 80'h10100000010000010010;
mem[728]  = 80'h00109400000208004500;
mem[729]  = 80'h0010002f5f3c0000fffd;
mem[730]  = 80'h0010da3cc0550102c000;
mem[731]  = 80'h00100001ffabffabffab;
mem[732]  = 80'h0010ffc3ce14fe5e7fc6;
mem[733]  = 80'h00107ba0dc160cccb9c9;
mem[734]  = 80'h0010d68fe024de22a32f;
mem[735]  = 80'h01112100000000000000;
mem[736]  = 80'h00000000000000000000;
mem[737]  = 80'h10100000010000010010;
mem[738]  = 80'h00109400000208004500;
mem[739]  = 80'h0010002f5f3d0000fffd;
mem[740]  = 80'h0010da3bc0550102c000;
mem[741]  = 80'h00100001ffabffabffab;
mem[742]  = 80'h0010ffc2bfcad2860604;
mem[743]  = 80'h0010c46b0e91e1396948;
mem[744]  = 80'h001087d683923e239513;
mem[745]  = 80'h01112100000000000000;
mem[746]  = 80'h00000000000000000000;
mem[747]  = 80'h00000000000000000000;
mem[748]  = 80'h00000000000000000000;
mem[749]  = 80'h10100000010000010010;
mem[750]  = 80'h00109400000208004500;
mem[751]  = 80'h0010002f5f3e0000fffd;
mem[752]  = 80'h0010da3ac0550102c000;
mem[753]  = 80'h00100001ffabffabffab;
mem[754]  = 80'h0010ffc12da8a7ee8c43;
mem[755]  = 80'h001004377919d72719cb;
mem[756]  = 80'h0010751a370683142473;
mem[757]  = 80'h0111c100000000000000;
mem[758]  = 80'h00000000000000000000;
mem[759]  = 80'h00000000000000000000;
mem[760]  = 80'h00000000000000000000;
mem[761]  = 80'h10100000010000010010;
mem[762]  = 80'h00109400000208004500;
mem[763]  = 80'h0010002f5f3f0000fffd;
mem[764]  = 80'h0010da39c0550102c000;
mem[765]  = 80'h00100001ffabffabffab;
mem[766]  = 80'h0010ffc05c768b36f581;
mem[767]  = 80'h0010bbfcab9e3ad2c9cd;
mem[768]  = 80'h001024c15b1436f98bcc;
mem[769]  = 80'h01116700000000000000;
mem[770]  = 80'h00000000000000000000;
mem[771]  = 80'h10100000010000010010;
mem[772]  = 80'h00109400000208004500;
mem[773]  = 80'h0010002f5f400000fffd;
mem[774]  = 80'h0010da38c0550102c000;
mem[775]  = 80'h00100001ffabffabffab;
mem[776]  = 80'h0010ffbfcbd386ed1e21;
mem[777]  = 80'h0010715ff320177b6e07;
mem[778]  = 80'h001043a410b750d62d19;
mem[779]  = 80'h01118000000000000000;
mem[780]  = 80'h00000000000000000000;
mem[781]  = 80'h00000000000000000000;
mem[782]  = 80'h00000000000000000000;
mem[783]  = 80'h10100000010000010010;
mem[784]  = 80'h00109400000208004500;
mem[785]  = 80'h0010002f5f410000fffd;
mem[786]  = 80'h0010da37c0550102c000;
mem[787]  = 80'h00100001ffabffabffab;
mem[788]  = 80'h0010ffbeba0daa3567e3;
mem[789]  = 80'h0010ce9421a7fa8ebd9e;
mem[790]  = 80'h0010122ef9827f1aacde;
mem[791]  = 80'h0111ed00000000000000;
mem[792]  = 80'h00000000000000000000;
mem[793]  = 80'h10100000010000010010;
mem[794]  = 80'h00109400000208004500;
mem[795]  = 80'h0010002f5f420000fffd;
mem[796]  = 80'h0010da36c0550102c000;
mem[797]  = 80'h00100001ffabffabffab;
mem[798]  = 80'h0010ffbd286fdf5deda4;
mem[799]  = 80'h00100ec8562fcc90cd15;
mem[800]  = 80'h0010e06be4c6463882f8;
mem[801]  = 80'h0111cc00000000000000;
mem[802]  = 80'h00000000000000000000;
mem[803]  = 80'h00000000000000000000;
mem[804]  = 80'h00000000000000000000;
mem[805]  = 80'h10100000010000010010;
mem[806]  = 80'h00109400000208004500;
mem[807]  = 80'h0010002f5f430000fffd;
mem[808]  = 80'h0010da35c0550102c000;
mem[809]  = 80'h00100001ffabffabffab;
mem[810]  = 80'h0010ffbc59b1f3859466;
mem[811]  = 80'h0010b10384a821651d1c;
mem[812]  = 80'h0010b1a0b6d7416681bf;
mem[813]  = 80'h0111eb00000000000000;
mem[814]  = 80'h00000000000000000000;
mem[815]  = 80'h10100000010000010010;
mem[816]  = 80'h00109400000208004500;
mem[817]  = 80'h0010002f5f440000fffd;
mem[818]  = 80'h0010da34c0550102c000;
mem[819]  = 80'h00100001ffabffabffab;
mem[820]  = 80'h0010ffbb7d75195480e9;
mem[821]  = 80'h001031bb6bb94d59fc67;
mem[822]  = 80'h001054314a2a623e745a;
mem[823]  = 80'h01111c00000000000000;
mem[824]  = 80'h00000000000000000000;
mem[825]  = 80'h00000000000000000000;
mem[826]  = 80'h00000000000000000000;
mem[827]  = 80'h00000000000000000000;
mem[828]  = 80'h10100000010000010010;
mem[829]  = 80'h00109400000208004500;
mem[830]  = 80'h0010002f5f450000fffd;
mem[831]  = 80'h0010da33c0550102c000;
mem[832]  = 80'h00100001ffabffabffab;
mem[833]  = 80'h0010ffba0cab358cf92b;
mem[834]  = 80'h00108e70b93ea0ac2c1e;
mem[835]  = 80'h001005f24176681352d0;
mem[836]  = 80'h01119500000000000000;
mem[837]  = 80'h10100000010000010010;
mem[838]  = 80'h00109400000208004500;
mem[839]  = 80'h0010002f5f460000fffd;
mem[840]  = 80'h0010da32c0550102c000;
mem[841]  = 80'h00100001ffabffabffab;
mem[842]  = 80'h0010ffb99ec940e4736c;
mem[843]  = 80'h00104e2cceb696b25c54;
mem[844]  = 80'h0010f79239af6b02ca51;
mem[845]  = 80'h0111b500000000000000;
mem[846]  = 80'h00000000000000000000;
mem[847]  = 80'h00000000000000000000;
mem[848]  = 80'h00000000000000000000;
mem[849]  = 80'h10100000010000010010;
mem[850]  = 80'h00109400000208004500;
mem[851]  = 80'h0010002f5f470000fffd;
mem[852]  = 80'h0010da31c0550102c000;
mem[853]  = 80'h00100001ffabffabffab;
mem[854]  = 80'h0010ffb8ef176c3c0aae;
mem[855]  = 80'h0010f1e71c317b478c1d;
mem[856]  = 80'h0010a654a77236615460;
mem[857]  = 80'h01111b00000000000000;
mem[858]  = 80'h10100000010000010010;
mem[859]  = 80'h00109400000208004500;
mem[860]  = 80'h0010002f5f480000fffd;
mem[861]  = 80'h0010da30c0550102c000;
mem[862]  = 80'h00100001ffabffabffab;
mem[863]  = 80'h0010ffb7d74095465a73;
mem[864]  = 80'h00104f5d10944ecb9ea3;
mem[865]  = 80'h00103cb1c13bed04127e;
mem[866]  = 80'h01115a00000000000000;
mem[867]  = 80'h00000000000000000000;
mem[868]  = 80'h00000000000000000000;
mem[869]  = 80'h00000000000000000000;
mem[870]  = 80'h10100000010000010010;
mem[871]  = 80'h00109400000208004500;
mem[872]  = 80'h0010002f5f490000fffd;
mem[873]  = 80'h0010da2fc0550102c000;
mem[874]  = 80'h00100001ffabffabffab;
mem[875]  = 80'h0010ffb6a69eb99e23b1;
mem[876]  = 80'h0010f096c213a33e4efa;
mem[877]  = 80'h00106d742c033dca842a;
mem[878]  = 80'h0111aa00000000000000;
mem[879]  = 80'h00000000000000000000;
mem[880]  = 80'h10100000010000010010;
mem[881]  = 80'h00109400000208004500;
mem[882]  = 80'h0010002f5f4a0000fffd;
mem[883]  = 80'h0010da2ec0550102c000;
mem[884]  = 80'h00100001ffabffabffab;
mem[885]  = 80'h0010ffb534fcccf6a9f6;
mem[886]  = 80'h001030cab59b95203fb1;
mem[887]  = 80'h00109f105518a43cf636;
mem[888]  = 80'h01118000000000000000;
mem[889]  = 80'h00000000000000000000;
mem[890]  = 80'h00000000000000000000;
mem[891]  = 80'h00000000000000000000;
mem[892]  = 80'h00000000000000000000;
mem[893]  = 80'h10100000010000010010;
mem[894]  = 80'h00109400000208004500;
mem[895]  = 80'h0010002f5f4b0000fffd;
mem[896]  = 80'h0010da2dc0550102c000;
mem[897]  = 80'h00100001ffabffabffab;
mem[898]  = 80'h0010ffb44522e02ed034;
mem[899]  = 80'h00108f01671c78d5eff8;
mem[900]  = 80'h0010ced6cb02119c436d;
mem[901]  = 80'h01110400000000000000;
mem[902]  = 80'h00000000000000000000;
mem[903]  = 80'h10100000010000010010;
mem[904]  = 80'h00109400000208004500;
mem[905]  = 80'h0010002f5f4c0000fffd;
mem[906]  = 80'h0010da2cc0550102c000;
mem[907]  = 80'h00100001ffabffabffab;
mem[908]  = 80'h0010ffb361e60affc4bb;
mem[909]  = 80'h00100fb9880d14e90ec0;
mem[910]  = 80'h00102b1fa81c3f14ca50;
mem[911]  = 80'h01118900000000000000;
mem[912]  = 80'h00000000000000000000;
mem[913]  = 80'h00000000000000000000;
mem[914]  = 80'h00000000000000000000;
mem[915]  = 80'h10100000010000010010;
mem[916]  = 80'h00109400000208004500;
mem[917]  = 80'h0010002f5f4d0000fffd;
mem[918]  = 80'h0010da2bc0550102c000;
mem[919]  = 80'h00100001ffabffabffab;
mem[920]  = 80'h0010ffb210382627bd79;
mem[921]  = 80'h0010b0725a8af91cdeb9;
mem[922]  = 80'h00107adca3c40a4b9c53;
mem[923]  = 80'h0111e900000000000000;
mem[924]  = 80'h00000000000000000000;
mem[925]  = 80'h10100000010000010010;
mem[926]  = 80'h00109400000208004500;
mem[927]  = 80'h0010002f5f4e0000fffd;
mem[928]  = 80'h0010da2ac0550102c000;
mem[929]  = 80'h00100001ffabffabffab;
mem[930]  = 80'h0010ffb1825a534f373e;
mem[931]  = 80'h0010702e2d02cf02ae32;
mem[932]  = 80'h00108899be6691c72489;
mem[933]  = 80'h0111f800000000000000;
mem[934]  = 80'h00000000000000000000;
mem[935]  = 80'h10100000010000010010;
mem[936]  = 80'h00109400000208004500;
mem[937]  = 80'h0010002f5f4f0000fffd;
mem[938]  = 80'h0010da29c0550102c000;
mem[939]  = 80'h00100001ffabffabffab;
mem[940]  = 80'h0010ffb0f3847f974efc;
mem[941]  = 80'h0010cfe5ff8522f77ebb;
mem[942]  = 80'h0010d94974ce7e2c75b0;
mem[943]  = 80'h01112e00000000000000;
mem[944]  = 80'h00000000000000000000;
mem[945]  = 80'h00000000000000000000;
mem[946]  = 80'h00000000000000000000;
mem[947]  = 80'h10100000010000010010;
mem[948]  = 80'h00109400000208004500;
mem[949]  = 80'h0010002f5f500000fffd;
mem[950]  = 80'h0010da28c0550102c000;
mem[951]  = 80'h00100001ffabffabffab;
mem[952]  = 80'h0010ffaff2f5a1bb9685;
mem[953]  = 80'h00100d5a3448a41a8b4f;
mem[954]  = 80'h0010bc4353c95319888a;
mem[955]  = 80'h01119f00000000000000;
mem[956]  = 80'h00000000000000000000;
mem[957]  = 80'h10100000010000010010;
mem[958]  = 80'h00109400000208004500;
mem[959]  = 80'h0010002f5f510000fffd;
mem[960]  = 80'h0010da27c0550102c000;
mem[961]  = 80'h00100001ffabffabffab;
mem[962]  = 80'h0010ffae832b8d63ef47;
mem[963]  = 80'h0010b291e6cf49ef5b56;
mem[964]  = 80'h0010ed8b724761744b83;
mem[965]  = 80'h01111700000000000000;
mem[966]  = 80'h00000000000000000000;
mem[967]  = 80'h00000000000000000000;
mem[968]  = 80'h00000000000000000000;
mem[969]  = 80'h10100000010000010010;
mem[970]  = 80'h00109400000208004500;
mem[971]  = 80'h0010002f5f520000fffd;
mem[972]  = 80'h0010da26c0550102c000;
mem[973]  = 80'h00100001ffabffabffab;
mem[974]  = 80'h0010ffad1149f80b6500;
mem[975]  = 80'h001072cd91477ff12bdc;
mem[976]  = 80'h00101ffd5e1d63e0b884;
mem[977]  = 80'h01115f00000000000000;
mem[978]  = 80'h00000000000000000000;
mem[979]  = 80'h10100000010000010010;
mem[980]  = 80'h00109400000208004500;
mem[981]  = 80'h0010002f5f530000fffd;
mem[982]  = 80'h0010da25c0550102c000;
mem[983]  = 80'h00100001ffabffabffab;
mem[984]  = 80'h0010ffac6097d4d31cc2;
mem[985]  = 80'h0010cd0643c092048455;
mem[986]  = 80'h00104ed9ad2b8a871482;
mem[987]  = 80'h0111b700000000000000;
mem[988]  = 80'h00000000000000000000;
mem[989]  = 80'h00000000000000000000;
mem[990]  = 80'h00000000000000000000;
mem[991]  = 80'h00000000000000000000;
mem[992]  = 80'h10100000010000010010;
mem[993]  = 80'h00109400000208004500;
mem[994]  = 80'h0010002f5f540000fffd;
mem[995]  = 80'h0010da24c0550102c000;
mem[996]  = 80'h00100001ffabffabffab;
mem[997]  = 80'h0010ffab44533e02084d;
mem[998]  = 80'h00104dbeacd1fe38652e;
mem[999]  = 80'h0010ab4851721a047a64;
mem[1000] = 80'h0111d800000000000000;
mem[1001] = 80'h10100000010000010010;
mem[1002] = 80'h00109400000208004500;
mem[1003] = 80'h0010002f5f550000fffd;
mem[1004] = 80'h0010da23c0550102c000;
mem[1005] = 80'h00100001ffabffabffab;
mem[1006] = 80'h0010ffaa358d12da718f;
mem[1007] = 80'h0010f2757e5613cdb557;
mem[1008] = 80'h0010fa8b5ae1b6759139;
mem[1009] = 80'h01112200000000000000;
mem[1010] = 80'h00000000000000000000;
mem[1011] = 80'h00000000000000000000;
mem[1012] = 80'h00000000000000000000;
mem[1013] = 80'h10100000010000010010;
mem[1014] = 80'h00109400000208004500;
mem[1015] = 80'h0010002f5f560000fffd;
mem[1016] = 80'h0010da22c0550102c000;
mem[1017] = 80'h00100001ffabffabffab;
mem[1018] = 80'h0010ffa9a7ef67b2fbc8;
mem[1019] = 80'h0010322909de25d3c59c;
mem[1020] = 80'h001008c38bb138b8f333;
mem[1021] = 80'h01111d00000000000000;
mem[1022] = 80'h00000000000000000000;
mem[1023] = 80'h10100000010000010010;
mem[1024] = 80'h00109400000208004500;
mem[1025] = 80'h0010002f5f570000fffd;
mem[1026] = 80'h0010da21c0550102c000;
mem[1027] = 80'h00100001ffabffabffab;
mem[1028] = 80'h0010ffa8d6314b6a820a;
mem[1029] = 80'h00108de2db59c82615d5;
mem[1030] = 80'h001059051573a64ff035;
mem[1031] = 80'h01117c00000000000000;
mem[1032] = 80'h00000000000000000000;
mem[1033] = 80'h00000000000000000000;
mem[1034] = 80'h00000000000000000000;
mem[1035] = 80'h10100000010000010010;
mem[1036] = 80'h00109400000208004500;
mem[1037] = 80'h0010002f5f580000fffd;
mem[1038] = 80'h0010da20c0550102c000;
mem[1039] = 80'h00100001ffabffabffab;
mem[1040] = 80'h0010ffa7ee66b210d2d7;
mem[1041] = 80'h00103358d7fcfdaa07ec;
mem[1042] = 80'h0010c3627cba3b29d7ae;
mem[1043] = 80'h0111d600000000000000;
mem[1044] = 80'h00000000000000000000;
mem[1045] = 80'h10100000010000010010;
mem[1046] = 80'h00109400000208004500;
mem[1047] = 80'h0010002f5f590000fffd;
mem[1048] = 80'h0010da1fc0550102c000;
mem[1049] = 80'h00100001ffabffabffab;
mem[1050] = 80'h0010ffa69fb89ec8ab15;
mem[1051] = 80'h00108c93057b105fd7ad;
mem[1052] = 80'h0010922d4b79be5c783f;
mem[1053] = 80'h01113e00000000000000;
mem[1054] = 80'h00000000000000000000;
mem[1055] = 80'h00000000000000000000;
mem[1056] = 80'h00000000000000000000;
mem[1057] = 80'h00000000000000000000;
mem[1058] = 80'h10100000010000010010;
mem[1059] = 80'h00109400000208004500;
mem[1060] = 80'h0010002f5f5a0000fffd;
mem[1061] = 80'h0010da1ec0550102c000;
mem[1062] = 80'h00100001ffabffabffab;
mem[1063] = 80'h0010ffa50ddaeba02152;
mem[1064] = 80'h00104ccf72f32641a77e;
mem[1065] = 80'h001060ef401bb6ba0ee1;
mem[1066] = 80'h01110500000000000000;
mem[1067] = 80'h10100000010000010010;
mem[1068] = 80'h00109400000208004500;
mem[1069] = 80'h0010002f5f5b0000fffd;
mem[1070] = 80'h0010da1dc0550102c000;
mem[1071] = 80'h00100001ffabffabffab;
mem[1072] = 80'h0010ffa47c04c7785890;
mem[1073] = 80'h0010f304a074cbb4773f;
mem[1074] = 80'h001031a0773fe48fcaba;
mem[1075] = 80'h01115400000000000000;
mem[1076] = 80'h00000000000000000000;
mem[1077] = 80'h00000000000000000000;
mem[1078] = 80'h00000000000000000000;
mem[1079] = 80'h10100000010000010010;
mem[1080] = 80'h00109400000208004500;
mem[1081] = 80'h0010002f5f5c0000fffd;
mem[1082] = 80'h0010da1cc0550102c000;
mem[1083] = 80'h00100001ffabffabffab;
mem[1084] = 80'h0010ffa358c02da94c1f;
mem[1085] = 80'h001073bc4f65a788978c;
mem[1086] = 80'h0010d4994603103b3d6d;
mem[1087] = 80'h01112300000000000000;
mem[1088] = 80'h00000000000000000000;
mem[1089] = 80'h10100000010000010010;
mem[1090] = 80'h00109400000208004500;
mem[1091] = 80'h0010002f5f5d0000fffd;
mem[1092] = 80'h0010da1bc0550102c000;
mem[1093] = 80'h00100001ffabffabffab;
mem[1094] = 80'h0010ffa2291e017135dd;
mem[1095] = 80'h0010cc779de24a7d47cd;
mem[1096] = 80'h001085d67175ab93c43d;
mem[1097] = 80'h01111b00000000000000;
mem[1098] = 80'h00000000000000000000;
mem[1099] = 80'h00000000000000000000;
mem[1100] = 80'h00000000000000000000;
mem[1101] = 80'h10100000010000010010;
mem[1102] = 80'h00109400000208004500;
mem[1103] = 80'h0010002f5f5e0000fffd;
mem[1104] = 80'h0010da1ac0550102c000;
mem[1105] = 80'h00100001ffabffabffab;
mem[1106] = 80'h0010ffa1bb7c7419bf9a;
mem[1107] = 80'h00100c2bea6a7c63377e;
mem[1108] = 80'h0010771f50969e031c3c;
mem[1109] = 80'h0111b000000000000000;
mem[1110] = 80'h00000000000000000000;
mem[1111] = 80'h00000000000000000000;
mem[1112] = 80'h00000000000000000000;
mem[1113] = 80'h10100000010000010010;
mem[1114] = 80'h00109400000208004500;
mem[1115] = 80'h0010002f5f5f0000fffd;
mem[1116] = 80'h0010da19c0550102c000;
mem[1117] = 80'h00100001ffabffabffab;
mem[1118] = 80'h0010ffa0caa258c1c658;
mem[1119] = 80'h0010b3e038ed9196e77e;
mem[1120] = 80'h0010266e9a50eff28ea4;
mem[1121] = 80'h01114600000000000000;
mem[1122] = 80'h00000000000000000000;
mem[1123] = 80'h10100000010000010010;
mem[1124] = 80'h00109400000208004500;
mem[1125] = 80'h0010002f5f600000fffd;
mem[1126] = 80'h0010da18c0550102c000;
mem[1127] = 80'h00100001ffabffabffab;
mem[1128] = 80'h0010ff9fb99fc8400f69;
mem[1129] = 80'h001089547df171b8dc97;
mem[1130] = 80'h0010bd382f482c41d142;
mem[1131] = 80'h0111ee00000000000000;
mem[1132] = 80'h00000000000000000000;
mem[1133] = 80'h00000000000000000000;
mem[1134] = 80'h00000000000000000000;
mem[1135] = 80'h10100000010000010010;
mem[1136] = 80'h00109400000208004500;
mem[1137] = 80'h0010002f5f610000fffd;
mem[1138] = 80'h0010da17c0550102c000;
mem[1139] = 80'h00100001ffabffabffab;
mem[1140] = 80'h0010ff9ec841e49876ab;
mem[1141] = 80'h0010369faf769c4d0c16;
mem[1142] = 80'h0010ec614c00152df0ee;
mem[1143] = 80'h0111eb00000000000000;
mem[1144] = 80'h00000000000000000000;
mem[1145] = 80'h10100000010000010010;
mem[1146] = 80'h00109400000208004500;
mem[1147] = 80'h0010002f5f620000fffd;
mem[1148] = 80'h0010da16c0550102c000;
mem[1149] = 80'h00100001ffabffabffab;
mem[1150] = 80'h0010ff9d5a2391f0fcec;
mem[1151] = 80'h0010f6c3d8feaa537c85;
mem[1152] = 80'h00101eae8b17763d0e9f;
mem[1153] = 80'h01113d00000000000000;
mem[1154] = 80'h00000000000000000000;
mem[1155] = 80'h00000000000000000000;
mem[1156] = 80'h00000000000000000000;
mem[1157] = 80'h10100000010000010010;
mem[1158] = 80'h00109400000208004500;
mem[1159] = 80'h0010002f5f630000fffd;
mem[1160] = 80'h0010da15c0550102c000;
mem[1161] = 80'h00100001ffabffabffab;
mem[1162] = 80'h0010ff9c2bfdbd28852e;
mem[1163] = 80'h001049080a7947a6ac84;
mem[1164] = 80'h00104fec70768988132a;
mem[1165] = 80'h01112c00000000000000;
mem[1166] = 80'h00000000000000000000;
mem[1167] = 80'h10100000010000010010;
mem[1168] = 80'h00109400000208004500;
mem[1169] = 80'h0010002f5f640000fffd;
mem[1170] = 80'h0010da14c0550102c000;
mem[1171] = 80'h00100001ffabffabffab;
mem[1172] = 80'h0010ff9b0f3957f991a1;
mem[1173] = 80'h0010c9b0e5682b9a4df7;
mem[1174] = 80'h0010aaf425f10dd45c06;
mem[1175] = 80'h0111ec00000000000000;
mem[1176] = 80'h00000000000000000000;
mem[1177] = 80'h00000000000000000000;
mem[1178] = 80'h00000000000000000000;
mem[1179] = 80'h00000000000000000000;
mem[1180] = 80'h10100000010000010010;
mem[1181] = 80'h00109400000208004500;
mem[1182] = 80'h0010002f5f650000fffd;
mem[1183] = 80'h0010da13c0550102c000;
mem[1184] = 80'h00100001ffabffabffab;
mem[1185] = 80'h0010ff9a7ee77b21e863;
mem[1186] = 80'h0010767b37efc66f9e75;
mem[1187] = 80'h0010fba14506c99299b7;
mem[1188] = 80'h0111c600000000000000;
mem[1189] = 80'h10100000010000010010;
mem[1190] = 80'h00109400000208004500;
mem[1191] = 80'h0010002f5f660000fffd;
mem[1192] = 80'h0010da12c0550102c000;
mem[1193] = 80'h00100001ffabffabffab;
mem[1194] = 80'h0010ff99ec850e496224;
mem[1195] = 80'h0010b6274067f071eec6;
mem[1196] = 80'h0010096864435f3fa834;
mem[1197] = 80'h0111da00000000000000;
mem[1198] = 80'h00000000000000000000;
mem[1199] = 80'h00000000000000000000;
mem[1200] = 80'h00000000000000000000;
mem[1201] = 80'h10100000010000010010;
mem[1202] = 80'h00109400000208004500;
mem[1203] = 80'h0010002f5f670000fffd;
mem[1204] = 80'h0010da11c0550102c000;
mem[1205] = 80'h00100001ffabffabffab;
mem[1206] = 80'h0010ff989d5b22911be6;
mem[1207] = 80'h001009ec92e01d843e87;
mem[1208] = 80'h0010582753957f25ffee;
mem[1209] = 80'h01111300000000000000;
mem[1210] = 80'h10100000010000010010;
mem[1211] = 80'h00109400000208004500;
mem[1212] = 80'h0010002f5f680000fffd;
mem[1213] = 80'h0010da10c0550102c000;
mem[1214] = 80'h00100001ffabffabffab;
mem[1215] = 80'h0010ff97a50cdbeb4b3b;
mem[1216] = 80'h0010b7569e4528082c31;
mem[1217] = 80'h0010c24b9c132b43f13e;
mem[1218] = 80'h0111c900000000000000;
mem[1219] = 80'h00000000000000000000;
mem[1220] = 80'h00000000000000000000;
mem[1221] = 80'h00000000000000000000;
mem[1222] = 80'h10100000010000010010;
mem[1223] = 80'h00109400000208004500;
mem[1224] = 80'h0010002f5f690000fffd;
mem[1225] = 80'h0010da0fc0550102c000;
mem[1226] = 80'h00100001ffabffabffab;
mem[1227] = 80'h0010ff96d4d2f73332f9;
mem[1228] = 80'h0010089d4cc2c5fdfc70;
mem[1229] = 80'h00109304ab96aa55b012;
mem[1230] = 80'h01119900000000000000;
mem[1231] = 80'h00000000000000000000;
mem[1232] = 80'h10100000010000010010;
mem[1233] = 80'h00109400000208004500;
mem[1234] = 80'h0010002f5f6a0000fffd;
mem[1235] = 80'h0010da0ec0550102c000;
mem[1236] = 80'h00100001ffabffabffab;
mem[1237] = 80'h0010ff9546b0825bb8be;
mem[1238] = 80'h0010c8c13b4af3e38c23;
mem[1239] = 80'h001061dd38af5f83e127;
mem[1240] = 80'h01115200000000000000;
mem[1241] = 80'h00000000000000000000;
mem[1242] = 80'h00000000000000000000;
mem[1243] = 80'h00000000000000000000;
mem[1244] = 80'h00000000000000000000;
mem[1245] = 80'h10100000010000010010;
mem[1246] = 80'h00109400000208004500;
mem[1247] = 80'h0010002f5f6b0000fffd;
mem[1248] = 80'h0010da0dc0550102c000;
mem[1249] = 80'h00100001ffabffabffab;
mem[1250] = 80'h0010ff94376eae83c17c;
mem[1251] = 80'h0010770ae9cd1e165c63;
mem[1252] = 80'h001030a13e0a0e4bd686;
mem[1253] = 80'h0111b400000000000000;
mem[1254] = 80'h00000000000000000000;
mem[1255] = 80'h10100000010000010010;
mem[1256] = 80'h00109400000208004500;
mem[1257] = 80'h0010002f5f6c0000fffd;
mem[1258] = 80'h0010da0cc0550102c000;
mem[1259] = 80'h00100001ffabffabffab;
mem[1260] = 80'h0010ff9313aa4452d5f3;
mem[1261] = 80'h0010f7b206dc722abd50;
mem[1262] = 80'h0010d5b4a7bd26b2fd0b;
mem[1263] = 80'h01111100000000000000;
mem[1264] = 80'h00000000000000000000;
mem[1265] = 80'h00000000000000000000;
mem[1266] = 80'h00000000000000000000;
mem[1267] = 80'h10100000010000010010;
mem[1268] = 80'h00109400000208004500;
mem[1269] = 80'h0010002f5f6d0000fffd;
mem[1270] = 80'h0010da0bc0550102c000;
mem[1271] = 80'h00100001ffabffabffab;
mem[1272] = 80'h0010ff926274688aac31;
mem[1273] = 80'h00104879d45b9fdf6d11;
mem[1274] = 80'h001084fb907b496fbc20;
mem[1275] = 80'h01114c00000000000000;
mem[1276] = 80'h00000000000000000000;
mem[1277] = 80'h10100000010000010010;
mem[1278] = 80'h00109400000208004500;
mem[1279] = 80'h0010002f5f6e0000fffd;
mem[1280] = 80'h0010da0ac0550102c000;
mem[1281] = 80'h00100001ffabffabffab;
mem[1282] = 80'h0010ff91f0161de22676;
mem[1283] = 80'h00108825a3d3a9c11da2;
mem[1284] = 80'h00107632b16fb01e9d0e;
mem[1285] = 80'h01112e00000000000000;
mem[1286] = 80'h00000000000000000000;
mem[1287] = 80'h10100000010000010010;
mem[1288] = 80'h00109400000208004500;
mem[1289] = 80'h0010002f5f6f0000fffd;
mem[1290] = 80'h0010da09c0550102c000;
mem[1291] = 80'h00100001ffabffabffab;
mem[1292] = 80'h0010ff9081c8313a5fb4;
mem[1293] = 80'h001037ee71544434cc23;
mem[1294] = 80'h0010275ce2c129758c40;
mem[1295] = 80'h01115200000000000000;
mem[1296] = 80'h00000000000000000000;
mem[1297] = 80'h00000000000000000000;
mem[1298] = 80'h00000000000000000000;
mem[1299] = 80'h10100000010000010010;
mem[1300] = 80'h00109400000208004500;
mem[1301] = 80'h0010002f5f700000fffd;
mem[1302] = 80'h0010da08c0550102c000;
mem[1303] = 80'h00100001ffabffabffab;
mem[1304] = 80'h0010ff8f80b9ef1687cd;
mem[1305] = 80'h0010f551ba99c2d939df;
mem[1306] = 80'h001042df6c4eacea5586;
mem[1307] = 80'h01116200000000000000;
mem[1308] = 80'h00000000000000000000;
mem[1309] = 80'h10100000010000010010;
mem[1310] = 80'h00109400000208004500;
mem[1311] = 80'h0010002f5f710000fffd;
mem[1312] = 80'h0010da07c0550102c000;
mem[1313] = 80'h00100001ffabffabffab;
mem[1314] = 80'h0010ff8ef167c3cefe0f;
mem[1315] = 80'h00104a9a681e2f2ce9d9;
mem[1316] = 80'h0010130400686d6c558b;
mem[1317] = 80'h01116000000000000000;
mem[1318] = 80'h00000000000000000000;
mem[1319] = 80'h00000000000000000000;
mem[1320] = 80'h00000000000000000000;
mem[1321] = 80'h10100000010000010010;
mem[1322] = 80'h00109400000208004500;
mem[1323] = 80'h0010002f5f720000fffd;
mem[1324] = 80'h0010da06c0550102c000;
mem[1325] = 80'h00100001ffabffabffab;
mem[1326] = 80'h0010ff8d6305b6a67448;
mem[1327] = 80'h00108ac61f9619329952;
mem[1328] = 80'h0010e1411d5b16c3b401;
mem[1329] = 80'h0111b900000000000000;
mem[1330] = 80'h00000000000000000000;
mem[1331] = 80'h10100000010000010010;
mem[1332] = 80'h00109400000208004500;
mem[1333] = 80'h0010002f5f730000fffd;
mem[1334] = 80'h0010da05c0550102c000;
mem[1335] = 80'h00100001ffabffabffab;
mem[1336] = 80'h0010ff8c12db9a7e0d8a;
mem[1337] = 80'h0010350dcd11f4c749cb;
mem[1338] = 80'h0010b092a44aaf647fe3;
mem[1339] = 80'h01119f00000000000000;
mem[1340] = 80'h00000000000000000000;
mem[1341] = 80'h00000000000000000000;
mem[1342] = 80'h00000000000000000000;
mem[1343] = 80'h00000000000000000000;
mem[1344] = 80'h10100000010000010010;
mem[1345] = 80'h00109400000208004500;
mem[1346] = 80'h0010002f5f740000fffd;
mem[1347] = 80'h0010da04c0550102c000;
mem[1348] = 80'h00100001ffabffabffab;
mem[1349] = 80'h0010ff8b361f70af1905;
mem[1350] = 80'h0010b5b5220098fba8b0;
mem[1351] = 80'h00105503583b79e85be7;
mem[1352] = 80'h01113200000000000000;
mem[1353] = 80'h10100000010000010010;
mem[1354] = 80'h00109400000208004500;
mem[1355] = 80'h0010002f5f750000fffd;
mem[1356] = 80'h0010da03c0550102c000;
mem[1357] = 80'h00100001ffabffabffab;
mem[1358] = 80'h0010ff8a47c15c7760c7;
mem[1359] = 80'h00100a7ef087750e78b9;
mem[1360] = 80'h001004c80ae002f20256;
mem[1361] = 80'h01114500000000000000;
mem[1362] = 80'h00000000000000000000;
mem[1363] = 80'h00000000000000000000;
mem[1364] = 80'h00000000000000000000;
mem[1365] = 80'h10100000010000010010;
mem[1366] = 80'h00109400000208004500;
mem[1367] = 80'h0010002f5f760000fffd;
mem[1368] = 80'h0010da02c0550102c000;
mem[1369] = 80'h00100001ffabffabffab;
mem[1370] = 80'h0010ff89d5a3291fea80;
mem[1371] = 80'h0010ca22870f43100832;
mem[1372] = 80'h0010f68d17306c99a752;
mem[1373] = 80'h01118400000000000000;
mem[1374] = 80'h00000000000000000000;
mem[1375] = 80'h10100000010000010010;
mem[1376] = 80'h00109400000208004500;
mem[1377] = 80'h0010002f5f770000fffd;
mem[1378] = 80'h0010da01c0550102c000;
mem[1379] = 80'h00100001ffabffabffab;
mem[1380] = 80'h0010ff88a47d05c79342;
mem[1381] = 80'h001075e95588aee5d84b;
mem[1382] = 80'h0010a74e1cfeabb68f2a;
mem[1383] = 80'h01119300000000000000;
mem[1384] = 80'h00000000000000000000;
mem[1385] = 80'h00000000000000000000;
mem[1386] = 80'h00000000000000000000;
mem[1387] = 80'h10100000010000010010;
mem[1388] = 80'h00109400000208004500;
mem[1389] = 80'h0010002f5f780000fffd;
mem[1390] = 80'h0010da00c0550102c000;
mem[1391] = 80'h00100001ffabffabffab;
mem[1392] = 80'h0010ff879c2afcbdc39f;
mem[1393] = 80'h0010cb53592d9b69cd74;
mem[1394] = 80'h00103d06438a95ae714c;
mem[1395] = 80'h0111ec00000000000000;
mem[1396] = 80'h00000000000000000000;
mem[1397] = 80'h10100000010000010010;
mem[1398] = 80'h00109400000208004500;
mem[1399] = 80'h0010002f5f790000fffd;
mem[1400] = 80'h0010d9ffc0550102c000;
mem[1401] = 80'h00100001ffabffabffab;
mem[1402] = 80'h0010ff86edf4d065ba5d;
mem[1403] = 80'h001074988baa769c1d3d;
mem[1404] = 80'h00106cc0dde3a8431d6d;
mem[1405] = 80'h01113100000000000000;
mem[1406] = 80'h00000000000000000000;
mem[1407] = 80'h00000000000000000000;
mem[1408] = 80'h00000000000000000000;
mem[1409] = 80'h00000000000000000000;
mem[1410] = 80'h10100000010000010010;
mem[1411] = 80'h00109400000208004500;
mem[1412] = 80'h0010002f5f7a0000fffd;
mem[1413] = 80'h0010d9fec0550102c000;
mem[1414] = 80'h00100001ffabffabffab;
mem[1415] = 80'h0010ff857f96a50d301a;
mem[1416] = 80'h0010b4c4fc2240826df6;
mem[1417] = 80'h00109e880cd3a03c3241;
mem[1418] = 80'h01116f00000000000000;
mem[1419] = 80'h10100000010000010010;
mem[1420] = 80'h00109400000208004500;
mem[1421] = 80'h0010002f5f7b0000fffd;
mem[1422] = 80'h0010d9fdc0550102c000;
mem[1423] = 80'h00100001ffabffabffab;
mem[1424] = 80'h0010ff840e4889d549d8;
mem[1425] = 80'h00100b0f2ea5ad77bdaf;
mem[1426] = 80'h0010cf4de15bc811badb;
mem[1427] = 80'h01111700000000000000;
mem[1428] = 80'h00000000000000000000;
mem[1429] = 80'h00000000000000000000;
mem[1430] = 80'h00000000000000000000;
mem[1431] = 80'h10100000010000010010;
mem[1432] = 80'h00109400000208004500;
mem[1433] = 80'h0010002f5f7c0000fffd;
mem[1434] = 80'h0010d9fcc0550102c000;
mem[1435] = 80'h00100001ffabffabffab;
mem[1436] = 80'h0010ff832a8c63045d57;
mem[1437] = 80'h00108bb7c1b4c14b5c14;
mem[1438] = 80'h00102aca49fe355df718;
mem[1439] = 80'h0111fc00000000000000;
mem[1440] = 80'h00000000000000000000;
mem[1441] = 80'h10100000010000010010;
mem[1442] = 80'h00109400000208004500;
mem[1443] = 80'h0010002f5f7d0000fffd;
mem[1444] = 80'h0010d9fbc0550102c000;
mem[1445] = 80'h00100001ffabffabffab;
mem[1446] = 80'h0010ff825b524fdc2495;
mem[1447] = 80'h0010347c13332cbe8c5d;
mem[1448] = 80'h00107b0cd7e1dcf0f3b9;
mem[1449] = 80'h01115f00000000000000;
mem[1450] = 80'h00000000000000000000;
mem[1451] = 80'h00000000000000000000;
mem[1452] = 80'h00000000000000000000;
mem[1453] = 80'h10100000010000010010;
mem[1454] = 80'h00109400000208004500;
mem[1455] = 80'h0010002f5f7e0000fffd;
mem[1456] = 80'h0010d9fac0550102c000;
mem[1457] = 80'h00100001ffabffabffab;
mem[1458] = 80'h0010ff81c9303ab4aed2;
mem[1459] = 80'h0010f42064bb1aa0fc95;
mem[1460] = 80'h0010891155a2febb2281;
mem[1461] = 80'h0111ca00000000000000;
mem[1462] = 80'h00000000000000000000;
mem[1463] = 80'h00000000000000000000;
mem[1464] = 80'h00000000000000000000;
mem[1465] = 80'h10100000010000010010;
mem[1466] = 80'h00109400000208004500;
mem[1467] = 80'h0010002f5f7f0000fffd;
mem[1468] = 80'h0010d9f9c0550102c000;
mem[1469] = 80'h00100001ffabffabffab;
mem[1470] = 80'h0010ff80b8ee166cd710;
mem[1471] = 80'h00104bebb63cf7552cec;
mem[1472] = 80'h0010d8d25ed6fb3aefb9;
mem[1473] = 80'h0111b600000000000000;
mem[1474] = 80'h00000000000000000000;
mem[1475] = 80'h10100000010000010010;
mem[1476] = 80'h00109400000208004500;
mem[1477] = 80'h0010002f5f800000fffd;
mem[1478] = 80'h0010d9f8c0550102c000;
mem[1479] = 80'h00100001ffabffabffab;
mem[1480] = 80'h0010ff7f97a40ddb0051;
mem[1481] = 80'h0010dead0741ac066314;
mem[1482] = 80'h001017030ea33fe81a2f;
mem[1483] = 80'h01110700000000000000;
mem[1484] = 80'h00000000000000000000;
mem[1485] = 80'h00000000000000000000;
mem[1486] = 80'h00000000000000000000;
mem[1487] = 80'h10100000010000010010;
mem[1488] = 80'h00109400000208004500;
mem[1489] = 80'h0010002f5f810000fffd;
mem[1490] = 80'h0010d9f7c0550102c000;
mem[1491] = 80'h00100001ffabffabffab;
mem[1492] = 80'h0010ff7ee67a21037993;
mem[1493] = 80'h00106166d5c641f3b29d;
mem[1494] = 80'h001046e4f4cd175daba6;
mem[1495] = 80'h0111ee00000000000000;
mem[1496] = 80'h00000000000000000000;
mem[1497] = 80'h10100000010000010010;
mem[1498] = 80'h00109400000208004500;
mem[1499] = 80'h0010002f5f820000fffd;
mem[1500] = 80'h0010d9f6c0550102c000;
mem[1501] = 80'h00100001ffabffabffab;
mem[1502] = 80'h0010ff7d7418546bf3d4;
mem[1503] = 80'h0010a13aa24e77edc216;
mem[1504] = 80'h0010b4a1e9fa27ee174e;
mem[1505] = 80'h0111b200000000000000;
mem[1506] = 80'h00000000000000000000;
mem[1507] = 80'h00000000000000000000;
mem[1508] = 80'h00000000000000000000;
mem[1509] = 80'h10100000010000010010;
mem[1510] = 80'h00109400000208004500;
mem[1511] = 80'h0010002f5f830000fffd;
mem[1512] = 80'h0010d9f5c0550102c000;
mem[1513] = 80'h00100001ffabffabffab;
mem[1514] = 80'h0010ff7c05c678b38a16;
mem[1515] = 80'h00101ef170c99a18120f;
mem[1516] = 80'h0010e569c8a70db033ce;
mem[1517] = 80'h0111cb00000000000000;
mem[1518] = 80'h00000000000000000000;
mem[1519] = 80'h10100000010000010010;
mem[1520] = 80'h00109400000208004500;
mem[1521] = 80'h0010002f5f840000fffd;
mem[1522] = 80'h0010d9f4c0550102c000;
mem[1523] = 80'h00100001ffabffabffab;
mem[1524] = 80'h0010ff7b210292629e99;
mem[1525] = 80'h00109e499fd8f624f375;
mem[1526] = 80'h001000cb05fe7f2ad547;
mem[1527] = 80'h0111e600000000000000;
mem[1528] = 80'h00000000000000000000;
mem[1529] = 80'h00000000000000000000;
mem[1530] = 80'h00000000000000000000;
mem[1531] = 80'h00000000000000000000;
mem[1532] = 80'h10100000010000010010;
mem[1533] = 80'h00109400000208004500;
mem[1534] = 80'h0010002f5f850000fffd;
mem[1535] = 80'h0010d9f3c0550102c000;
mem[1536] = 80'h00100001ffabffabffab;
mem[1537] = 80'h0010ff7a50dcbebae75b;
mem[1538] = 80'h001021824d5f1bd123fc;
mem[1539] = 80'h0010511bcfc8398e60e6;
mem[1540] = 80'h01114800000000000000;
mem[1541] = 80'h10100000010000010010;
mem[1542] = 80'h00109400000208004500;
mem[1543] = 80'h0010002f5f860000fffd;
mem[1544] = 80'h0010d9f2c0550102c000;
mem[1545] = 80'h00100001ffabffabffab;
mem[1546] = 80'h0010ff79c2becbd26d1c;
mem[1547] = 80'h0010e1de3ad72dcf5377;
mem[1548] = 80'h0010a35ed27cf00d5dc1;
mem[1549] = 80'h0111c000000000000000;
mem[1550] = 80'h00000000000000000000;
mem[1551] = 80'h00000000000000000000;
mem[1552] = 80'h00000000000000000000;
mem[1553] = 80'h10100000010000010010;
mem[1554] = 80'h00109400000208004500;
mem[1555] = 80'h0010002f5f870000fffd;
mem[1556] = 80'h0010d9f1c0550102c000;
mem[1557] = 80'h00100001ffabffabffab;
mem[1558] = 80'h0010ff78b360e70a14de;
mem[1559] = 80'h00105e15e850c03a830e;
mem[1560] = 80'h0010f29dd9effa36e879;
mem[1561] = 80'h01113d00000000000000;
mem[1562] = 80'h10100000010000010010;
mem[1563] = 80'h00109400000208004500;
mem[1564] = 80'h0010002f5f880000fffd;
mem[1565] = 80'h0010d9f0c0550102c000;
mem[1566] = 80'h00100001ffabffabffab;
mem[1567] = 80'h0010ff778b371e704403;
mem[1568] = 80'h0010e0afe4f5f5b691b0;
mem[1569] = 80'h00106878bf579d088117;
mem[1570] = 80'h0111b300000000000000;
mem[1571] = 80'h00000000000000000000;
mem[1572] = 80'h00000000000000000000;
mem[1573] = 80'h00000000000000000000;
mem[1574] = 80'h10100000010000010010;
mem[1575] = 80'h00109400000208004500;
mem[1576] = 80'h0010002f5f890000fffd;
mem[1577] = 80'h0010d9efc0550102c000;
mem[1578] = 80'h00100001ffabffabffab;
mem[1579] = 80'h0010ff76fae932a83dc1;
mem[1580] = 80'h00105f643672184341f9;
mem[1581] = 80'h001039be216549294015;
mem[1582] = 80'h0111f900000000000000;
mem[1583] = 80'h00000000000000000000;
mem[1584] = 80'h10100000010000010010;
mem[1585] = 80'h00109400000208004500;
mem[1586] = 80'h0010002f5f8a0000fffd;
mem[1587] = 80'h0010d9eec0550102c000;
mem[1588] = 80'h00100001ffabffabffab;
mem[1589] = 80'h0010ff75688b47c0b786;
mem[1590] = 80'h00109f3841fa2e5d32b5;
mem[1591] = 80'h0010cb2daf44dbf45fd2;
mem[1592] = 80'h01114000000000000000;
mem[1593] = 80'h00000000000000000000;
mem[1594] = 80'h00000000000000000000;
mem[1595] = 80'h00000000000000000000;
mem[1596] = 80'h00000000000000000000;
mem[1597] = 80'h10100000010000010010;
mem[1598] = 80'h00109400000208004500;
mem[1599] = 80'h0010002f5f8b0000fffd;
mem[1600] = 80'h0010d9edc0550102c000;
mem[1601] = 80'h00100001ffabffabffab;
mem[1602] = 80'h0010ff7419556b18ce44;
mem[1603] = 80'h001020f3937dc3a8e2f4;
mem[1604] = 80'h00109a6298681fb8273c;
mem[1605] = 80'h0111c000000000000000;
mem[1606] = 80'h00000000000000000000;
mem[1607] = 80'h10100000010000010010;
mem[1608] = 80'h00109400000208004500;
mem[1609] = 80'h0010002f5f8c0000fffd;
mem[1610] = 80'h0010d9ecc0550102c000;
mem[1611] = 80'h00100001ffabffabffab;
mem[1612] = 80'h0010ff733d9181c9dacb;
mem[1613] = 80'h0010a04b7c6caf9403d7;
mem[1614] = 80'h00107f7472cda3b350f3;
mem[1615] = 80'h0111ad00000000000000;
mem[1616] = 80'h00000000000000000000;
mem[1617] = 80'h00000000000000000000;
mem[1618] = 80'h00000000000000000000;
mem[1619] = 80'h10100000010000010010;
mem[1620] = 80'h00109400000208004500;
mem[1621] = 80'h0010002f5f8d0000fffd;
mem[1622] = 80'h0010d9ebc0550102c000;
mem[1623] = 80'h00100001ffabffabffab;
mem[1624] = 80'h0010ff724c4fad11a309;
mem[1625] = 80'h00101f80aeeb4261d396;
mem[1626] = 80'h00102e3b45840bf9c2c3;
mem[1627] = 80'h01114900000000000000;
mem[1628] = 80'h00000000000000000000;
mem[1629] = 80'h10100000010000010010;
mem[1630] = 80'h00109400000208004500;
mem[1631] = 80'h0010002f5f8e0000fffd;
mem[1632] = 80'h0010d9eac0550102c000;
mem[1633] = 80'h00100001ffabffabffab;
mem[1634] = 80'h0010ff71de2dd879294e;
mem[1635] = 80'h0010dfdcd963747fa3d5;
mem[1636] = 80'h0010dce1a520cc844d1a;
mem[1637] = 80'h0111c900000000000000;
mem[1638] = 80'h00000000000000000000;
mem[1639] = 80'h10100000010000010010;
mem[1640] = 80'h00109400000208004500;
mem[1641] = 80'h0010002f5f8f0000fffd;
mem[1642] = 80'h0010d9e9c0550102c000;
mem[1643] = 80'h00100001ffabffabffab;
mem[1644] = 80'h0010ff70aff3f4a1508c;
mem[1645] = 80'h001060170be4998a7394;
mem[1646] = 80'h00108dae92a471b1caf3;
mem[1647] = 80'h01110600000000000000;
mem[1648] = 80'h00000000000000000000;
mem[1649] = 80'h00000000000000000000;
mem[1650] = 80'h00000000000000000000;
mem[1651] = 80'h10100000010000010010;
mem[1652] = 80'h00109400000208004500;
mem[1653] = 80'h0010002f5f900000fffd;
mem[1654] = 80'h0010d9e8c0550102c000;
mem[1655] = 80'h00100001ffabffabffab;
mem[1656] = 80'h0010ff6fae822a8d88f5;
mem[1657] = 80'h0010a2a8c0291f678658;
mem[1658] = 80'h0010e82889d023abe1b6;
mem[1659] = 80'h01111100000000000000;
mem[1660] = 80'h00000000000000000000;
mem[1661] = 80'h10100000010000010010;
mem[1662] = 80'h00109400000208004500;
mem[1663] = 80'h0010002f5f910000fffd;
mem[1664] = 80'h0010d9e7c0550102c000;
mem[1665] = 80'h00100001ffabffabffab;
mem[1666] = 80'h0010ff6edf5c0655f137;
mem[1667] = 80'h00101d6312aef2925658;
mem[1668] = 80'h0010b9594351b3cf91eb;
mem[1669] = 80'h0111c700000000000000;
mem[1670] = 80'h00000000000000000000;
mem[1671] = 80'h00000000000000000000;
mem[1672] = 80'h00000000000000000000;
mem[1673] = 80'h10100000010000010010;
mem[1674] = 80'h00109400000208004500;
mem[1675] = 80'h0010002f5f920000fffd;
mem[1676] = 80'h0010d9e6c0550102c000;
mem[1677] = 80'h00100001ffabffabffab;
mem[1678] = 80'h0010ff6d4d3e733d7b70;
mem[1679] = 80'h0010dd3f6526c48c26db;
mem[1680] = 80'h00104b95f742533d0393;
mem[1681] = 80'h01114600000000000000;
mem[1682] = 80'h00000000000000000000;
mem[1683] = 80'h10100000010000010010;
mem[1684] = 80'h00109400000208004500;
mem[1685] = 80'h0010002f5f930000fffd;
mem[1686] = 80'h0010d9e5c0550102c000;
mem[1687] = 80'h00100001ffabffabffab;
mem[1688] = 80'h0010ff6c3ce05fe502b2;
mem[1689] = 80'h001062f4b7a12979f75a;
mem[1690] = 80'h00101afba4b665f119e0;
mem[1691] = 80'h01113c00000000000000;
mem[1692] = 80'h00000000000000000000;
mem[1693] = 80'h00000000000000000000;
mem[1694] = 80'h00000000000000000000;
mem[1695] = 80'h00000000000000000000;
mem[1696] = 80'h10100000010000010010;
mem[1697] = 80'h00109400000208004500;
mem[1698] = 80'h0010002f5f940000fffd;
mem[1699] = 80'h0010d9e4c0550102c000;
mem[1700] = 80'h00100001ffabffabffab;
mem[1701] = 80'h0010ff6b1824b534163d;
mem[1702] = 80'h0010e24c58b045451639;
mem[1703] = 80'h0010ffe082a2035c7770;
mem[1704] = 80'h0111af00000000000000;
mem[1705] = 80'h10100000010000010010;
mem[1706] = 80'h00109400000208004500;
mem[1707] = 80'h0010002f5f950000fffd;
mem[1708] = 80'h0010d9e3c0550102c000;
mem[1709] = 80'h00100001ffabffabffab;
mem[1710] = 80'h0010ff6a69fa99ec6fff;
mem[1711] = 80'h00105d878a37a8b0c638;
mem[1712] = 80'h0010aea279640ddada69;
mem[1713] = 80'h0111ad00000000000000;
mem[1714] = 80'h00000000000000000000;
mem[1715] = 80'h00000000000000000000;
mem[1716] = 80'h00000000000000000000;
mem[1717] = 80'h10100000010000010010;
mem[1718] = 80'h00109400000208004500;
mem[1719] = 80'h0010002f5f960000fffd;
mem[1720] = 80'h0010d9e2c0550102c000;
mem[1721] = 80'h00100001ffabffabffab;
mem[1722] = 80'h0010ff69fb98ec84e5b8;
mem[1723] = 80'h00109ddbfdbf9eaeb6bb;
mem[1724] = 80'h00105c6ecd4b17d52a8a;
mem[1725] = 80'h01110200000000000000;
mem[1726] = 80'h00000000000000000000;
mem[1727] = 80'h10100000010000010010;
mem[1728] = 80'h00109400000208004500;
mem[1729] = 80'h0010002f5f970000fffd;
mem[1730] = 80'h0010d9e1c0550102c000;
mem[1731] = 80'h00100001ffabffabffab;
mem[1732] = 80'h0010ff688a46c05c9c7a;
mem[1733] = 80'h001022102f38735b6639;
mem[1734] = 80'h00100d62fd39e3a39f17;
mem[1735] = 80'h01119b00000000000000;
mem[1736] = 80'h00000000000000000000;
mem[1737] = 80'h00000000000000000000;
mem[1738] = 80'h00000000000000000000;
mem[1739] = 80'h10100000010000010010;
mem[1740] = 80'h00109400000208004500;
mem[1741] = 80'h0010002f5f980000fffd;
mem[1742] = 80'h0010d9e0c0550102c000;
mem[1743] = 80'h00100001ffabffabffab;
mem[1744] = 80'h0010ff67b2113926cca7;
mem[1745] = 80'h00109caa239d46d774ff;
mem[1746] = 80'h001097066b93c94196b0;
mem[1747] = 80'h01116200000000000000;
mem[1748] = 80'h00000000000000000000;
mem[1749] = 80'h10100000010000010010;
mem[1750] = 80'h00109400000208004500;
mem[1751] = 80'h0010002f5f990000fffd;
mem[1752] = 80'h0010d9dfc0550102c000;
mem[1753] = 80'h00100001ffabffabffab;
mem[1754] = 80'h0010ff66c3cf15feb565;
mem[1755] = 80'h00102361f11aab22a4be;
mem[1756] = 80'h0010c6495cbee931b060;
mem[1757] = 80'h0111ec00000000000000;
mem[1758] = 80'h00000000000000000000;
mem[1759] = 80'h00000000000000000000;
mem[1760] = 80'h00000000000000000000;
mem[1761] = 80'h00000000000000000000;
mem[1762] = 80'h10100000010000010010;
mem[1763] = 80'h00109400000208004500;
mem[1764] = 80'h0010002f5f9a0000fffd;
mem[1765] = 80'h0010d9dec0550102c000;
mem[1766] = 80'h00100001ffabffabffab;
mem[1767] = 80'h0010ff6551ad60963f22;
mem[1768] = 80'h0010e33d86929d3cd47d;
mem[1769] = 80'h001034882421da7fcb73;
mem[1770] = 80'h01118000000000000000;
mem[1771] = 80'h10100000010000010010;
mem[1772] = 80'h00109400000208004500;
mem[1773] = 80'h0010002f5f9b0000fffd;
mem[1774] = 80'h0010d9ddc0550102c000;
mem[1775] = 80'h00100001ffabffabffab;
mem[1776] = 80'h0010ff6420734c4e46e0;
mem[1777] = 80'h00105cf6541570c9043c;
mem[1778] = 80'h001065c71321adab3ac4;
mem[1779] = 80'h01116b00000000000000;
mem[1780] = 80'h00000000000000000000;
mem[1781] = 80'h00000000000000000000;
mem[1782] = 80'h00000000000000000000;
mem[1783] = 80'h10100000010000010010;
mem[1784] = 80'h00109400000208004500;
mem[1785] = 80'h0010002f5f9c0000fffd;
mem[1786] = 80'h0010d9dcc0550102c000;
mem[1787] = 80'h00100001ffabffabffab;
mem[1788] = 80'h0010ff6304b7a69f526f;
mem[1789] = 80'h0010dc4ebb041cf5ea9f;
mem[1790] = 80'h001080e65007927496b9;
mem[1791] = 80'h01113100000000000000;
mem[1792] = 80'h00000000000000000000;
mem[1793] = 80'h10100000010000010010;
mem[1794] = 80'h00109400000208004500;
mem[1795] = 80'h0010002f5f9d0000fffd;
mem[1796] = 80'h0010d9dbc0550102c000;
mem[1797] = 80'h00100001ffabffabffab;
mem[1798] = 80'h0010ff6275698a472bad;
mem[1799] = 80'h001063856983f1003adf;
mem[1800] = 80'h0010d19a56bbb30f214d;
mem[1801] = 80'h01112400000000000000;
mem[1802] = 80'h00000000000000000000;
mem[1803] = 80'h00000000000000000000;
mem[1804] = 80'h00000000000000000000;
mem[1805] = 80'h10100000010000010010;
mem[1806] = 80'h00109400000208004500;
mem[1807] = 80'h0010002f5f9e0000fffd;
mem[1808] = 80'h0010d9dac0550102c000;
mem[1809] = 80'h00100001ffabffabffab;
mem[1810] = 80'h0010ff61e70bff2fa1ea;
mem[1811] = 80'h0010a3d91e0bc71e4a1c;
mem[1812] = 80'h0010235b2efd52ef9779;
mem[1813] = 80'h01117000000000000000;
mem[1814] = 80'h00000000000000000000;
mem[1815] = 80'h00000000000000000000;
mem[1816] = 80'h00000000000000000000;
mem[1817] = 80'h10100000010000010010;
mem[1818] = 80'h00109400000208004500;
mem[1819] = 80'h0010002f5f9f0000fffd;
mem[1820] = 80'h0010d9d9c0550102c000;
mem[1821] = 80'h00100001ffabffabffab;
mem[1822] = 80'h0010ff6096d5d3f7d828;
mem[1823] = 80'h00101c12cc8c2aeb9a5d;
mem[1824] = 80'h0010721419ad83b23dc0;
mem[1825] = 80'h01111e00000000000000;
mem[1826] = 80'h00000000000000000000;
mem[1827] = 80'h10100000010000010010;
mem[1828] = 80'h00109400000208004500;
mem[1829] = 80'h0010002f5fa00000fffd;
mem[1830] = 80'h0010d9d8c0550102c000;
mem[1831] = 80'h00100001ffabffabffab;
mem[1832] = 80'h0010ff5fe5e843761119;
mem[1833] = 80'h001026a68990cac5a184;
mem[1834] = 80'h0010e947395f866693cc;
mem[1835] = 80'h0111a800000000000000;
mem[1836] = 80'h00000000000000000000;
mem[1837] = 80'h00000000000000000000;
mem[1838] = 80'h00000000000000000000;
mem[1839] = 80'h10100000010000010010;
mem[1840] = 80'h00109400000208004500;
mem[1841] = 80'h0010002f5fa10000fffd;
mem[1842] = 80'h0010d9d7c0550102c000;
mem[1843] = 80'h00100001ffabffabffab;
mem[1844] = 80'h0010ff5e94366fae68db;
mem[1845] = 80'h0010996d5b1727307105;
mem[1846] = 80'h0010b81e5a07f44338ac;
mem[1847] = 80'h01110600000000000000;
mem[1848] = 80'h00000000000000000000;
mem[1849] = 80'h10100000010000010010;
mem[1850] = 80'h00109400000208004500;
mem[1851] = 80'h0010002f5fa20000fffd;
mem[1852] = 80'h0010d9d6c0550102c000;
mem[1853] = 80'h00100001ffabffabffab;
mem[1854] = 80'h0010ff5d06541ac6e29c;
mem[1855] = 80'h001059312c9f112e0186;
mem[1856] = 80'h00104ad2ee942a512f36;
mem[1857] = 80'h01117d00000000000000;
mem[1858] = 80'h00000000000000000000;
mem[1859] = 80'h00000000000000000000;
mem[1860] = 80'h00000000000000000000;
mem[1861] = 80'h10100000010000010010;
mem[1862] = 80'h00109400000208004500;
mem[1863] = 80'h0010002f5fa30000fffd;
mem[1864] = 80'h0010d9d5c0550102c000;
mem[1865] = 80'h00100001ffabffabffab;
mem[1866] = 80'h0010ff5c778a361e9b5e;
mem[1867] = 80'h0010e6fafe18fcdbd180;
mem[1868] = 80'h00101b09822266e9b383;
mem[1869] = 80'h0111d500000000000000;
mem[1870] = 80'h00000000000000000000;
mem[1871] = 80'h10100000010000010010;
mem[1872] = 80'h00109400000208004500;
mem[1873] = 80'h0010002f5fa40000fffd;
mem[1874] = 80'h0010d9d4c0550102c000;
mem[1875] = 80'h00100001ffabffabffab;
mem[1876] = 80'h0010ff5b534edccf8fd1;
mem[1877] = 80'h00106642110990e730fb;
mem[1878] = 80'h0010fe987eed895b9cc4;
mem[1879] = 80'h01115d00000000000000;
mem[1880] = 80'h00000000000000000000;
mem[1881] = 80'h00000000000000000000;
mem[1882] = 80'h00000000000000000000;
mem[1883] = 80'h00000000000000000000;
mem[1884] = 80'h10100000010000010010;
mem[1885] = 80'h00109400000208004500;
mem[1886] = 80'h0010002f5fa50000fffd;
mem[1887] = 80'h0010d9d3c0550102c000;
mem[1888] = 80'h00100001ffabffabffab;
mem[1889] = 80'h0010ff5a2290f017f613;
mem[1890] = 80'h0010d989c38e7d12e162;
mem[1891] = 80'h0010af7cf7de5436c2fb;
mem[1892] = 80'h01114100000000000000;
mem[1893] = 80'h10100000010000010010;
mem[1894] = 80'h00109400000208004500;
mem[1895] = 80'h0010002f5fa60000fffd;
mem[1896] = 80'h0010d9d2c0550102c000;
mem[1897] = 80'h00100001ffabffabffab;
mem[1898] = 80'h0010ff59b0f2857f7c54;
mem[1899] = 80'h001019d5b4064b0c91e9;
mem[1900] = 80'h00105d39ead45a902b9a;
mem[1901] = 80'h0111b600000000000000;
mem[1902] = 80'h00000000000000000000;
mem[1903] = 80'h00000000000000000000;
mem[1904] = 80'h00000000000000000000;
mem[1905] = 80'h10100000010000010010;
mem[1906] = 80'h00109400000208004500;
mem[1907] = 80'h0010002f5fa70000fffd;
mem[1908] = 80'h0010d9d1c0550102c000;
mem[1909] = 80'h00100001ffabffabffab;
mem[1910] = 80'h0010ff58c12ca9a70596;
mem[1911] = 80'h0010a61e6681a6f941e0;
mem[1912] = 80'h00100cf2b8d0d45ef50c;
mem[1913] = 80'h01113200000000000000;
mem[1914] = 80'h10100000010000010010;
mem[1915] = 80'h00109400000208004500;
mem[1916] = 80'h0010002f5fa80000fffd;
mem[1917] = 80'h0010d9d0c0550102c000;
mem[1918] = 80'h00100001ffabffabffab;
mem[1919] = 80'h0010ff57f97b50dd554b;
mem[1920] = 80'h001018a46a249375531e;
mem[1921] = 80'h0010961a128d4efda8e0;
mem[1922] = 80'h01113900000000000000;
mem[1923] = 80'h00000000000000000000;
mem[1924] = 80'h00000000000000000000;
mem[1925] = 80'h00000000000000000000;
mem[1926] = 80'h10100000010000010010;
mem[1927] = 80'h00109400000208004500;
mem[1928] = 80'h0010002f5fa90000fffd;
mem[1929] = 80'h0010d9cfc0550102c000;
mem[1930] = 80'h00100001ffabffabffab;
mem[1931] = 80'h0010ff5688a57c052c89;
mem[1932] = 80'h0010a76fb8a37e808367;
mem[1933] = 80'h0010c7d919a08b34ca74;
mem[1934] = 80'h01111c00000000000000;
mem[1935] = 80'h00000000000000000000;
mem[1936] = 80'h10100000010000010010;
mem[1937] = 80'h00109400000208004500;
mem[1938] = 80'h0010002f5faa0000fffd;
mem[1939] = 80'h0010d9cec0550102c000;
mem[1940] = 80'h00100001ffabffabffab;
mem[1941] = 80'h0010ff551ac7096da6ce;
mem[1942] = 80'h00106733cf2b489ef32d;
mem[1943] = 80'h001035b961c32b45e600;
mem[1944] = 80'h01116d00000000000000;
mem[1945] = 80'h00000000000000000000;
mem[1946] = 80'h00000000000000000000;
mem[1947] = 80'h00000000000000000000;
mem[1948] = 80'h00000000000000000000;
mem[1949] = 80'h10100000010000010010;
mem[1950] = 80'h00109400000208004500;
mem[1951] = 80'h0010002f5fab0000fffd;
mem[1952] = 80'h0010d9cdc0550102c000;
mem[1953] = 80'h00100001ffabffabffab;
mem[1954] = 80'h0010ff546b1925b5df0c;
mem[1955] = 80'h0010d8f81daca56b2364;
mem[1956] = 80'h0010647fffdb6c57a2de;
mem[1957] = 80'h01118800000000000000;
mem[1958] = 80'h00000000000000000000;
mem[1959] = 80'h10100000010000010010;
mem[1960] = 80'h00109400000208004500;
mem[1961] = 80'h0010002f5fac0000fffd;
mem[1962] = 80'h0010d9ccc0550102c000;
mem[1963] = 80'h00100001ffabffabffab;
mem[1964] = 80'h0010ff534fddcf64cb83;
mem[1965] = 80'h00105840f2bdc957c25f;
mem[1966] = 80'h001081e3cf4ced73ab76;
mem[1967] = 80'h0111bd00000000000000;
mem[1968] = 80'h00000000000000000000;
mem[1969] = 80'h00000000000000000000;
mem[1970] = 80'h00000000000000000000;
mem[1971] = 80'h10100000010000010010;
mem[1972] = 80'h00109400000208004500;
mem[1973] = 80'h0010002f5fad0000fffd;
mem[1974] = 80'h0010d9cbc0550102c000;
mem[1975] = 80'h00100001ffabffabffab;
mem[1976] = 80'h0010ff523e03e3bcb241;
mem[1977] = 80'h0010e78b203a24a21206;
mem[1978] = 80'h0010d0262216fb6f800f;
mem[1979] = 80'h0111f900000000000000;
mem[1980] = 80'h00000000000000000000;
mem[1981] = 80'h10100000010000010010;
mem[1982] = 80'h00109400000208004500;
mem[1983] = 80'h0010002f5fae0000fffd;
mem[1984] = 80'h0010d9cac0550102c000;
mem[1985] = 80'h00100001ffabffabffab;
mem[1986] = 80'h0010ff51ac6196d43806;
mem[1987] = 80'h001027d757b212bc614d;
mem[1988] = 80'h0010222c3bb333f44a88;
mem[1989] = 80'h0111b100000000000000;
mem[1990] = 80'h00000000000000000000;
mem[1991] = 80'h10100000010000010010;
mem[1992] = 80'h00109400000208004500;
mem[1993] = 80'h0010002f5faf0000fffd;
mem[1994] = 80'h0010d9c9c0550102c000;
mem[1995] = 80'h00100001ffabffabffab;
mem[1996] = 80'h0010ff50ddbfba0c41c4;
mem[1997] = 80'h0010981c8535ff49b104;
mem[1998] = 80'h001073eaa5933f052ac7;
mem[1999] = 80'h0111a200000000000000;
mem[2000] = 80'h00000000000000000000;
mem[2001] = 80'h00000000000000000000;
mem[2002] = 80'h00000000000000000000;
mem[2003] = 80'h10100000010000010010;
mem[2004] = 80'h00109400000208004500;
mem[2005] = 80'h0010002f5fb00000fffd;
mem[2006] = 80'h0010d9c8c0550102c000;
mem[2007] = 80'h00100001ffabffabffab;
mem[2008] = 80'h0010ff4fdcce642099bd;
mem[2009] = 80'h00105aa34ef879a444b3;
mem[2010] = 80'h001016b81d5889fca555;
mem[2011] = 80'h01116200000000000000;
mem[2012] = 80'h00000000000000000000;
mem[2013] = 80'h10100000010000010010;
mem[2014] = 80'h00109400000208004500;
mem[2015] = 80'h0010002f5fb10000fffd;
mem[2016] = 80'h0010d9c7c0550102c000;
mem[2017] = 80'h00100001ffabffabffab;
mem[2018] = 80'h0010ff4ead1048f8e07f;
mem[2019] = 80'h0010e5689c7f945194ca;
mem[2020] = 80'h0010477b16a920090209;
mem[2021] = 80'h0111cf00000000000000;
mem[2022] = 80'h00000000000000000000;
mem[2023] = 80'h00000000000000000000;
mem[2024] = 80'h00000000000000000000;
mem[2025] = 80'h10100000010000010010;
mem[2026] = 80'h00109400000208004500;
mem[2027] = 80'h0010002f5fb20000fffd;
mem[2028] = 80'h0010d9c6c0550102c000;
mem[2029] = 80'h00100001ffabffabffab;
mem[2030] = 80'h0010ff4d3f723d906a38;
mem[2031] = 80'h00102534ebf7a24fe441;
mem[2032] = 80'h0010b53e0b7bc0c76b3b;
mem[2033] = 80'h01113600000000000000;
mem[2034] = 80'h00000000000000000000;
mem[2035] = 80'h10100000010000010010;
mem[2036] = 80'h00109400000208004500;
mem[2037] = 80'h0010002f5fb30000fffd;
mem[2038] = 80'h0010d9c5c0550102c000;
mem[2039] = 80'h00100001ffabffabffab;
mem[2040] = 80'h0010ff4c4eac114813fa;
mem[2041] = 80'h00109aff39704fba34c8;
mem[2042] = 80'h0010e4eec1e38c8dfe9b;
mem[2043] = 80'h01117000000000000000;
mem[2044] = 80'h00000000000000000000;
mem[2045] = 80'h00000000000000000000;
mem[2046] = 80'h00000000000000000000;
mem[2047] = 80'h00000000000000000000;
mem[2048] = 80'h10100000010000010010;
mem[2049] = 80'h00109400000208004500;
mem[2050] = 80'h0010002f5fb40000fffd;
mem[2051] = 80'h0010d9c4c0550102c000;
mem[2052] = 80'h00100001ffabffabffab;
mem[2053] = 80'h0010ff4b6a68fb990775;
mem[2054] = 80'h00101a47d6612386d5b3;
mem[2055] = 80'h0010017f3ddb695b4ff4;
mem[2056] = 80'h01114300000000000000;
mem[2057] = 80'h10100000010000010010;
mem[2058] = 80'h00109400000208004500;
mem[2059] = 80'h0010002f5fb50000fffd;
mem[2060] = 80'h0010d9c3c0550102c000;
mem[2061] = 80'h00100001ffabffabffab;
mem[2062] = 80'h0010ff4a1bb6d7417eb7;
mem[2063] = 80'h0010a58c04e6ce7305aa;
mem[2064] = 80'h001050b71cbea2875db6;
mem[2065] = 80'h0111c200000000000000;
mem[2066] = 80'h00000000000000000000;
mem[2067] = 80'h00000000000000000000;
mem[2068] = 80'h00000000000000000000;
mem[2069] = 80'h10100000010000010010;
mem[2070] = 80'h00109400000208004500;
mem[2071] = 80'h0010002f5fb60000fffd;
mem[2072] = 80'h0010d9c2c0550102c000;
mem[2073] = 80'h00100001ffabffabffab;
mem[2074] = 80'h0010ff4989d4a229f4f0;
mem[2075] = 80'h001065d0736ef86d7520;
mem[2076] = 80'h0010a2c13038c5d7b1e4;
mem[2077] = 80'h01119a00000000000000;
mem[2078] = 80'h00000000000000000000;
mem[2079] = 80'h10100000010000010010;
mem[2080] = 80'h00109400000208004500;
mem[2081] = 80'h0010002f5fb70000fffd;
mem[2082] = 80'h0010d9c1c0550102c000;
mem[2083] = 80'h00100001ffabffabffab;
mem[2084] = 80'h0010ff48f80a8ef18d32;
mem[2085] = 80'h0010da1ba1e91598a4a9;
mem[2086] = 80'h0010f326ca19f8fa5ea1;
mem[2087] = 80'h01112100000000000000;
mem[2088] = 80'h00000000000000000000;
mem[2089] = 80'h00000000000000000000;
mem[2090] = 80'h00000000000000000000;
mem[2091] = 80'h10100000010000010010;
mem[2092] = 80'h00109400000208004500;
mem[2093] = 80'h0010002f5fb80000fffd;
mem[2094] = 80'h0010d9c0c0550102c000;
mem[2095] = 80'h00100001ffabffabffab;
mem[2096] = 80'h0010ff47c05d778bddef;
mem[2097] = 80'h001064a1ad4c2014b657;
mem[2098] = 80'h001069ce60b7375c14dd;
mem[2099] = 80'h01110e00000000000000;
mem[2100] = 80'h00000000000000000000;
mem[2101] = 80'h10100000010000010010;
mem[2102] = 80'h00109400000208004500;
mem[2103] = 80'h0010002f5fb90000fffd;
mem[2104] = 80'h0010d9bfc0550102c000;
mem[2105] = 80'h00100001ffabffabffab;
mem[2106] = 80'h0010ff46b1835b53a42d;
mem[2107] = 80'h0010db6a7fcbcde1662e;
mem[2108] = 80'h0010380d6b611c97c6a7;
mem[2109] = 80'h0111b100000000000000;
mem[2110] = 80'h00000000000000000000;
mem[2111] = 80'h00000000000000000000;
mem[2112] = 80'h00000000000000000000;
mem[2113] = 80'h00000000000000000000;
mem[2114] = 80'h10100000010000010010;
mem[2115] = 80'h00109400000208004500;
mem[2116] = 80'h0010002f5fba0000fffd;
mem[2117] = 80'h0010d9bec0550102c000;
mem[2118] = 80'h00100001ffabffabffab;
mem[2119] = 80'h0010ff4523e12e3b2e6a;
mem[2120] = 80'h00101b360843fbff16e5;
mem[2121] = 80'h0010ca45ba8fc4add3e3;
mem[2122] = 80'h01117600000000000000;
mem[2123] = 80'h10100000010000010010;
mem[2124] = 80'h00109400000208004500;
mem[2125] = 80'h0010002f5fbb0000fffd;
mem[2126] = 80'h0010d9bdc0550102c000;
mem[2127] = 80'h00100001ffabffabffab;
mem[2128] = 80'h0010ff44523f02e357a8;
mem[2129] = 80'h0010a4fddac4160ac6ac;
mem[2130] = 80'h00109b8324f436d8e8e6;
mem[2131] = 80'h01116600000000000000;
mem[2132] = 80'h00000000000000000000;
mem[2133] = 80'h00000000000000000000;
mem[2134] = 80'h00000000000000000000;
mem[2135] = 80'h10100000010000010010;
mem[2136] = 80'h00109400000208004500;
mem[2137] = 80'h0010002f5fbc0000fffd;
mem[2138] = 80'h0010d9bcc0550102c000;
mem[2139] = 80'h00100001ffabffabffab;
mem[2140] = 80'h0010ff4376fbe8324327;
mem[2141] = 80'h0010244535d57a362710;
mem[2142] = 80'h00107e9d1b68c87749b9;
mem[2143] = 80'h01113f00000000000000;
mem[2144] = 80'h00000000000000000000;
mem[2145] = 80'h10100000010000010010;
mem[2146] = 80'h00109400000208004500;
mem[2147] = 80'h0010002f5fbd0000fffd;
mem[2148] = 80'h0010d9bbc0550102c000;
mem[2149] = 80'h00100001ffabffabffab;
mem[2150] = 80'h0010ff420725c4ea3ae5;
mem[2151] = 80'h00109b8ee75297c3f751;
mem[2152] = 80'h00102fd22cff8aca38ed;
mem[2153] = 80'h01118400000000000000;
mem[2154] = 80'h00000000000000000000;
mem[2155] = 80'h00000000000000000000;
mem[2156] = 80'h00000000000000000000;
mem[2157] = 80'h10100000010000010010;
mem[2158] = 80'h00109400000208004500;
mem[2159] = 80'h0010002f5fbe0000fffd;
mem[2160] = 80'h0010d9bac0550102c000;
mem[2161] = 80'h00100001ffabffabffab;
mem[2162] = 80'h0010ff419547b182b0a2;
mem[2163] = 80'h00105bd290daa1dd8782;
mem[2164] = 80'h0010dd102733ee38f2b3;
mem[2165] = 80'h0111cb00000000000000;
mem[2166] = 80'h00000000000000000000;
mem[2167] = 80'h00000000000000000000;
mem[2168] = 80'h00000000000000000000;
mem[2169] = 80'h10100000010000010010;
mem[2170] = 80'h00109400000208004500;
mem[2171] = 80'h0010002f5fbf0000fffd;
mem[2172] = 80'h0010d9b9c0550102c000;
mem[2173] = 80'h00100001ffabffabffab;
mem[2174] = 80'h0010ff40e4999d5ac960;
mem[2175] = 80'h0010e419425d4c2857c3;
mem[2176] = 80'h00108c5f10a84df0460f;
mem[2177] = 80'h01113300000000000000;
mem[2178] = 80'h00000000000000000000;
mem[2179] = 80'h10100000010000010010;
mem[2180] = 80'h00109400000208004500;
mem[2181] = 80'h0010002f5fc00000fffd;
mem[2182] = 80'h0010d9b8c0550102c000;
mem[2183] = 80'h00100001ffabffabffab;
mem[2184] = 80'h0010ff3f733c908122c0;
mem[2185] = 80'h00102eba1ae36181f7c1;
mem[2186] = 80'h0010eb2036411524179a;
mem[2187] = 80'h01115800000000000000;
mem[2188] = 80'h00000000000000000000;
mem[2189] = 80'h00000000000000000000;
mem[2190] = 80'h00000000000000000000;
mem[2191] = 80'h10100000010000010010;
mem[2192] = 80'h00109400000208004500;
mem[2193] = 80'h0010002f5fc10000fffd;
mem[2194] = 80'h0010d9b7c0550102c000;
mem[2195] = 80'h00100001ffabffabffab;
mem[2196] = 80'h0010ff3e02e2bc595b02;
mem[2197] = 80'h00109171c8648c742780;
mem[2198] = 80'h0010ba6f01491c7ad9b9;
mem[2199] = 80'h01118400000000000000;
mem[2200] = 80'h00000000000000000000;
mem[2201] = 80'h10100000010000010010;
mem[2202] = 80'h00109400000208004500;
mem[2203] = 80'h0010002f5fc20000fffd;
mem[2204] = 80'h0010d9b6c0550102c000;
mem[2205] = 80'h00100001ffabffabffab;
mem[2206] = 80'h0010ff3d9080c931d145;
mem[2207] = 80'h0010512dbfecba6a5733;
mem[2208] = 80'h001048a6206c497a10aa;
mem[2209] = 80'h0111ff00000000000000;
mem[2210] = 80'h00000000000000000000;
mem[2211] = 80'h00000000000000000000;
mem[2212] = 80'h00000000000000000000;
mem[2213] = 80'h10100000010000010010;
mem[2214] = 80'h00109400000208004500;
mem[2215] = 80'h0010002f5fc30000fffd;
mem[2216] = 80'h0010d9b5c0550102c000;
mem[2217] = 80'h00100001ffabffabffab;
mem[2218] = 80'h0010ff3ce15ee5e9a887;
mem[2219] = 80'h0010eee66d6b579f8733;
mem[2220] = 80'h001019d7eaf650b97955;
mem[2221] = 80'h01115c00000000000000;
mem[2222] = 80'h00000000000000000000;
mem[2223] = 80'h10100000010000010010;
mem[2224] = 80'h00109400000208004500;
mem[2225] = 80'h0010002f5fc40000fffd;
mem[2226] = 80'h0010d9b4c0550102c000;
mem[2227] = 80'h00100001ffabffabffab;
mem[2228] = 80'h0010ff3bc59a0f38bc08;
mem[2229] = 80'h00106e5e827a3ba36640;
mem[2230] = 80'h0010fccfbf5c200f5a83;
mem[2231] = 80'h01110600000000000000;
mem[2232] = 80'h00000000000000000000;
mem[2233] = 80'h00000000000000000000;
mem[2234] = 80'h00000000000000000000;
mem[2235] = 80'h00000000000000000000;
mem[2236] = 80'h10100000010000010010;
mem[2237] = 80'h00109400000208004500;
mem[2238] = 80'h0010002f5fc50000fffd;
mem[2239] = 80'h0010d9b3c0550102c000;
mem[2240] = 80'h00100001ffabffabffab;
mem[2241] = 80'h0010ff3ab44423e0c5ca;
mem[2242] = 80'h0010d19550fdd656b6c1;
mem[2243] = 80'h0010ad96dc9328fbc493;
mem[2244] = 80'h01115600000000000000;
mem[2245] = 80'h10100000010000010010;
mem[2246] = 80'h00109400000208004500;
mem[2247] = 80'h0010002f5fc60000fffd;
mem[2248] = 80'h0010d9b2c0550102c000;
mem[2249] = 80'h00100001ffabffabffab;
mem[2250] = 80'h0010ff39262656884f8d;
mem[2251] = 80'h001011c92775e048c652;
mem[2252] = 80'h00105f591b57d95f5ef6;
mem[2253] = 80'h01113400000000000000;
mem[2254] = 80'h00000000000000000000;
mem[2255] = 80'h00000000000000000000;
mem[2256] = 80'h00000000000000000000;
mem[2257] = 80'h10100000010000010010;
mem[2258] = 80'h00109400000208004500;
mem[2259] = 80'h0010002f5fc70000fffd;
mem[2260] = 80'h0010d9b1c0550102c000;
mem[2261] = 80'h00100001ffabffabffab;
mem[2262] = 80'h0010ff3857f87a50364f;
mem[2263] = 80'h0010ae02f5f20dbd1653;
mem[2264] = 80'h00100e1be00e41ea0b0a;
mem[2265] = 80'h0111e100000000000000;
mem[2266] = 80'h10100000010000010010;
mem[2267] = 80'h00109400000208004500;
mem[2268] = 80'h0010002f5fc80000fffd;
mem[2269] = 80'h0010d9b0c0550102c000;
mem[2270] = 80'h00100001ffabffabffab;
mem[2271] = 80'h0010ff376faf832a6692;
mem[2272] = 80'h001010b8f957383104a5;
mem[2273] = 80'h0010947ae3fae75d30e7;
mem[2274] = 80'h01111000000000000000;
mem[2275] = 80'h00000000000000000000;
mem[2276] = 80'h00000000000000000000;
mem[2277] = 80'h00000000000000000000;
mem[2278] = 80'h10100000010000010010;
mem[2279] = 80'h00109400000208004500;
mem[2280] = 80'h0010002f5fc90000fffd;
mem[2281] = 80'h0010d9afc0550102c000;
mem[2282] = 80'h00100001ffabffabffab;
mem[2283] = 80'h0010ff361e71aff21f50;
mem[2284] = 80'h0010af732bd0d5c4d527;
mem[2285] = 80'h0010c541e3a2e3c61efd;
mem[2286] = 80'h01111d00000000000000;
mem[2287] = 80'h00000000000000000000;
mem[2288] = 80'h10100000010000010010;
mem[2289] = 80'h00109400000208004500;
mem[2290] = 80'h0010002f5fca0000fffd;
mem[2291] = 80'h0010d9aec0550102c000;
mem[2292] = 80'h00100001ffabffabffab;
mem[2293] = 80'h0010ff358c13da9a9517;
mem[2294] = 80'h00106f2f5c58e3daa594;
mem[2295] = 80'h00103788c284b5bfd5ca;
mem[2296] = 80'h0111d400000000000000;
mem[2297] = 80'h00000000000000000000;
mem[2298] = 80'h00000000000000000000;
mem[2299] = 80'h00000000000000000000;
mem[2300] = 80'h00000000000000000000;
mem[2301] = 80'h10100000010000010010;
mem[2302] = 80'h00109400000208004500;
mem[2303] = 80'h0010002f5fcb0000fffd;
mem[2304] = 80'h0010d9adc0550102c000;
mem[2305] = 80'h00100001ffabffabffab;
mem[2306] = 80'h0010ff34fdcdf642ecd5;
mem[2307] = 80'h0010d0e48edf0e2f75d5;
mem[2308] = 80'h001066c7f553df6a1b02;
mem[2309] = 80'h01119200000000000000;
mem[2310] = 80'h00000000000000000000;
mem[2311] = 80'h10100000010000010010;
mem[2312] = 80'h00109400000208004500;
mem[2313] = 80'h0010002f5fcc0000fffd;
mem[2314] = 80'h0010d9acc0550102c000;
mem[2315] = 80'h00100001ffabffabffab;
mem[2316] = 80'h0010ff33d9091c93f85a;
mem[2317] = 80'h0010505c61ce621394e6;
mem[2318] = 80'h001083d26cdd7898230c;
mem[2319] = 80'h01114400000000000000;
mem[2320] = 80'h00000000000000000000;
mem[2321] = 80'h00000000000000000000;
mem[2322] = 80'h00000000000000000000;
mem[2323] = 80'h10100000010000010010;
mem[2324] = 80'h00109400000208004500;
mem[2325] = 80'h0010002f5fcd0000fffd;
mem[2326] = 80'h0010d9abc0550102c000;
mem[2327] = 80'h00100001ffabffabffab;
mem[2328] = 80'h0010ff32a8d7304b8198;
mem[2329] = 80'h0010ef97b3498fe644a7;
mem[2330] = 80'h0010d29d5b05005dd8b5;
mem[2331] = 80'h01114e00000000000000;
mem[2332] = 80'h00000000000000000000;
mem[2333] = 80'h10100000010000010010;
mem[2334] = 80'h00109400000208004500;
mem[2335] = 80'h0010002f5fce0000fffd;
mem[2336] = 80'h0010d9aac0550102c000;
mem[2337] = 80'h00100001ffabffabffab;
mem[2338] = 80'h0010ff313ab545230bdf;
mem[2339] = 80'h00102fcbc4c1b9f834f4;
mem[2340] = 80'h00102044c858a8610acb;
mem[2341] = 80'h01119100000000000000;
mem[2342] = 80'h00000000000000000000;
mem[2343] = 80'h10100000010000010010;
mem[2344] = 80'h00109400000208004500;
mem[2345] = 80'h0010002f5fcf0000fffd;
mem[2346] = 80'h0010d9a9c0550102c000;
mem[2347] = 80'h00100001ffabffabffab;
mem[2348] = 80'h0010ff304b6b69fb721d;
mem[2349] = 80'h001090001646540de4b4;
mem[2350] = 80'h00107138ce09ba3a096f;
mem[2351] = 80'h0111e800000000000000;
mem[2352] = 80'h00000000000000000000;
mem[2353] = 80'h00000000000000000000;
mem[2354] = 80'h00000000000000000000;
mem[2355] = 80'h10100000010000010010;
mem[2356] = 80'h00109400000208004500;
mem[2357] = 80'h0010002f5fd00000fffd;
mem[2358] = 80'h0010d9a8c0550102c000;
mem[2359] = 80'h00100001ffabffabffab;
mem[2360] = 80'h0010ff2f4a1ab7d7aa64;
mem[2361] = 80'h001052bfdd8bd2e01108;
mem[2362] = 80'h001014b68c8f9e07453d;
mem[2363] = 80'h0111cd00000000000000;
mem[2364] = 80'h00000000000000000000;
mem[2365] = 80'h10100000010000010010;
mem[2366] = 80'h00109400000208004500;
mem[2367] = 80'h0010002f5fd10000fffd;
mem[2368] = 80'h0010d9a7c0550102c000;
mem[2369] = 80'h00100001ffabffabffab;
mem[2370] = 80'h0010ff2e3bc49b0fd3a6;
mem[2371] = 80'h0010ed740f0c3f15c149;
mem[2372] = 80'h001045f9bb7d57de4029;
mem[2373] = 80'h01116400000000000000;
mem[2374] = 80'h00000000000000000000;
mem[2375] = 80'h00000000000000000000;
mem[2376] = 80'h00000000000000000000;
mem[2377] = 80'h10100000010000010010;
mem[2378] = 80'h00109400000208004500;
mem[2379] = 80'h0010002f5fd20000fffd;
mem[2380] = 80'h0010d9a6c0550102c000;
mem[2381] = 80'h00100001ffabffabffab;
mem[2382] = 80'h0010ff2da9a6ee6759e1;
mem[2383] = 80'h00102d287884090bb1fa;
mem[2384] = 80'h0010b7309aff5ba04acb;
mem[2385] = 80'h0111ec00000000000000;
mem[2386] = 80'h00000000000000000000;
mem[2387] = 80'h10100000010000010010;
mem[2388] = 80'h00109400000208004500;
mem[2389] = 80'h0010002f5fd30000fffd;
mem[2390] = 80'h0010d9a5c0550102c000;
mem[2391] = 80'h00100001ffabffabffab;
mem[2392] = 80'h0010ff2cd878c2bf2023;
mem[2393] = 80'h001092e3aa03e4fe627b;
mem[2394] = 80'h0010e630a9e5307ef92e;
mem[2395] = 80'h01114700000000000000;
mem[2396] = 80'h00000000000000000000;
mem[2397] = 80'h00000000000000000000;
mem[2398] = 80'h00000000000000000000;
mem[2399] = 80'h00000000000000000000;
mem[2400] = 80'h10100000010000010010;
mem[2401] = 80'h00109400000208004500;
mem[2402] = 80'h0010002f5fd40000fffd;
mem[2403] = 80'h0010d9a4c0550102c000;
mem[2404] = 80'h00100001ffabffabffab;
mem[2405] = 80'h0010ff2bfcbc286e34ac;
mem[2406] = 80'h0010125b451288c28308;
mem[2407] = 80'h00100328fc9c43ae1de4;
mem[2408] = 80'h01112e00000000000000;
mem[2409] = 80'h10100000010000010010;
mem[2410] = 80'h00109400000208004500;
mem[2411] = 80'h0010002f5fd50000fffd;
mem[2412] = 80'h0010d9a3c0550102c000;
mem[2413] = 80'h00100001ffabffabffab;
mem[2414] = 80'h0010ff2a8d6204b64d6e;
mem[2415] = 80'h0010ad9097956537530e;
mem[2416] = 80'h001052f390ef3f26ca55;
mem[2417] = 80'h01112e00000000000000;
mem[2418] = 80'h00000000000000000000;
mem[2419] = 80'h00000000000000000000;
mem[2420] = 80'h00000000000000000000;
mem[2421] = 80'h10100000010000010010;
mem[2422] = 80'h00109400000208004500;
mem[2423] = 80'h0010002f5fd60000fffd;
mem[2424] = 80'h0010d9a2c0550102c000;
mem[2425] = 80'h00100001ffabffabffab;
mem[2426] = 80'h0010ff291f0071dec729;
mem[2427] = 80'h00106dcce01d53292385;
mem[2428] = 80'h0010a0b68d7eb5683754;
mem[2429] = 80'h0111a100000000000000;
mem[2430] = 80'h00000000000000000000;
mem[2431] = 80'h10100000010000010010;
mem[2432] = 80'h00109400000208004500;
mem[2433] = 80'h0010002f5fd70000fffd;
mem[2434] = 80'h0010d9a1c0550102c000;
mem[2435] = 80'h00100001ffabffabffab;
mem[2436] = 80'h0010ff286ede5d06beeb;
mem[2437] = 80'h0010d207329abedcf31c;
mem[2438] = 80'h0010f1653405992918c1;
mem[2439] = 80'h01119800000000000000;
mem[2440] = 80'h00000000000000000000;
mem[2441] = 80'h00000000000000000000;
mem[2442] = 80'h00000000000000000000;
mem[2443] = 80'h10100000010000010010;
mem[2444] = 80'h00109400000208004500;
mem[2445] = 80'h0010002f5fd80000fffd;
mem[2446] = 80'h0010d9a0c0550102c000;
mem[2447] = 80'h00100001ffabffabffab;
mem[2448] = 80'h0010ff275689a47cee36;
mem[2449] = 80'h00106cbd3e3f8b50e1e2;
mem[2450] = 80'h00106b8d9eddf43b4e00;
mem[2451] = 80'h0111f600000000000000;
mem[2452] = 80'h00000000000000000000;
mem[2453] = 80'h10100000010000010010;
mem[2454] = 80'h00109400000208004500;
mem[2455] = 80'h0010002f5fd90000fffd;
mem[2456] = 80'h0010d99fc0550102c000;
mem[2457] = 80'h00100001ffabffabffab;
mem[2458] = 80'h0010ff26275788a497f4;
mem[2459] = 80'h0010d376ecb866a531eb;
mem[2460] = 80'h00103a46cce258357706;
mem[2461] = 80'h01112b00000000000000;
mem[2462] = 80'h00000000000000000000;
mem[2463] = 80'h00000000000000000000;
mem[2464] = 80'h00000000000000000000;
mem[2465] = 80'h00000000000000000000;
mem[2466] = 80'h10100000010000010010;
mem[2467] = 80'h00109400000208004500;
mem[2468] = 80'h0010002f5fda0000fffd;
mem[2469] = 80'h0010d99ec0550102c000;
mem[2470] = 80'h00100001ffabffabffab;
mem[2471] = 80'h0010ff25b535fdcc1db3;
mem[2472] = 80'h0010132a9b3050bb4160;
mem[2473] = 80'h0010c803d1aa55aee221;
mem[2474] = 80'h01118700000000000000;
mem[2475] = 80'h10100000010000010010;
mem[2476] = 80'h00109400000208004500;
mem[2477] = 80'h0010002f5fdb0000fffd;
mem[2478] = 80'h0010d99dc0550102c000;
mem[2479] = 80'h00100001ffabffabffab;
mem[2480] = 80'h0010ff24c4ebd1146471;
mem[2481] = 80'h0010ace149b7bd4e9119;
mem[2482] = 80'h001099c0daa74cdfb1e5;
mem[2483] = 80'h01111100000000000000;
mem[2484] = 80'h00000000000000000000;
mem[2485] = 80'h00000000000000000000;
mem[2486] = 80'h00000000000000000000;
mem[2487] = 80'h10100000010000010010;
mem[2488] = 80'h00109400000208004500;
mem[2489] = 80'h0010002f5fdc0000fffd;
mem[2490] = 80'h0010d99cc0550102c000;
mem[2491] = 80'h00100001ffabffabffab;
mem[2492] = 80'h0010ff23e02f3bc570fe;
mem[2493] = 80'h00102c59a6a6d17271a3;
mem[2494] = 80'h00107c43738f6d1ba1e5;
mem[2495] = 80'h01111800000000000000;
mem[2496] = 80'h00000000000000000000;
mem[2497] = 80'h10100000010000010010;
mem[2498] = 80'h00109400000208004500;
mem[2499] = 80'h0010002f5fdd0000fffd;
mem[2500] = 80'h0010d99bc0550102c000;
mem[2501] = 80'h00100001ffabffabffab;
mem[2502] = 80'h0010ff2291f1171d093c;
mem[2503] = 80'h0010939274213c87a1ea;
mem[2504] = 80'h00102d85ede74c050085;
mem[2505] = 80'h01114e00000000000000;
mem[2506] = 80'h00000000000000000000;
mem[2507] = 80'h00000000000000000000;
mem[2508] = 80'h00000000000000000000;
mem[2509] = 80'h10100000010000010010;
mem[2510] = 80'h00109400000208004500;
mem[2511] = 80'h0010002f5fde0000fffd;
mem[2512] = 80'h0010d99ac0550102c000;
mem[2513] = 80'h00100001ffabffabffab;
mem[2514] = 80'h0010ff2103936275837b;
mem[2515] = 80'h001053ce03a90a99d121;
mem[2516] = 80'h0010dfcd3c5ac7e61b35;
mem[2517] = 80'h0111ea00000000000000;
mem[2518] = 80'h00000000000000000000;
mem[2519] = 80'h00000000000000000000;
mem[2520] = 80'h00000000000000000000;
mem[2521] = 80'h10100000010000010010;
mem[2522] = 80'h00109400000208004500;
mem[2523] = 80'h0010002f5fdf0000fffd;
mem[2524] = 80'h0010d999c0550102c000;
mem[2525] = 80'h00100001ffabffabffab;
mem[2526] = 80'h0010ff20724d4eadfab9;
mem[2527] = 80'h0010ec05d12ee76c0178;
mem[2528] = 80'h00108e08d1083f1a2d77;
mem[2529] = 80'h01111900000000000000;
mem[2530] = 80'h00000000000000000000;
mem[2531] = 80'h10100000010000010010;
mem[2532] = 80'h00109400000208004500;
mem[2533] = 80'h0010002f5fe00000fffd;
mem[2534] = 80'h0010d998c0550102c000;
mem[2535] = 80'h00100001ffabffabffab;
mem[2536] = 80'h0010ff1f0170de2c3388;
mem[2537] = 80'h0010d6b1943207423a59;
mem[2538] = 80'h001015c1997a91c96104;
mem[2539] = 80'h0111b800000000000000;
mem[2540] = 80'h00000000000000000000;
mem[2541] = 80'h00000000000000000000;
mem[2542] = 80'h00000000000000000000;
mem[2543] = 80'h10100000010000010010;
mem[2544] = 80'h00109400000208004500;
mem[2545] = 80'h0010002f5fe10000fffd;
mem[2546] = 80'h0010d997c0550102c000;
mem[2547] = 80'h00100001ffabffabffab;
mem[2548] = 80'h0010ff1e70aef2f44a4a;
mem[2549] = 80'h0010697a46b5eab7ea10;
mem[2550] = 80'h0010440707f481a9253e;
mem[2551] = 80'h0111c700000000000000;
mem[2552] = 80'h00000000000000000000;
mem[2553] = 80'h10100000010000010010;
mem[2554] = 80'h00109400000208004500;
mem[2555] = 80'h0010002f5fe20000fffd;
mem[2556] = 80'h0010d996c0550102c000;
mem[2557] = 80'h00100001ffabffabffab;
mem[2558] = 80'h0010ff1de2cc879cc00d;
mem[2559] = 80'h0010a926313ddca99ad8;
mem[2560] = 80'h0010b61a856a48407448;
mem[2561] = 80'h01115100000000000000;
mem[2562] = 80'h00000000000000000000;
mem[2563] = 80'h00000000000000000000;
mem[2564] = 80'h00000000000000000000;
mem[2565] = 80'h10100000010000010010;
mem[2566] = 80'h00109400000208004500;
mem[2567] = 80'h0010002f5fe30000fffd;
mem[2568] = 80'h0010d995c0550102c000;
mem[2569] = 80'h00100001ffabffabffab;
mem[2570] = 80'h0010ff1c9312ab44b9cf;
mem[2571] = 80'h001016ede3ba315c4aa1;
mem[2572] = 80'h0010e7d98e3d1b613ad1;
mem[2573] = 80'h01111100000000000000;
mem[2574] = 80'h00000000000000000000;
mem[2575] = 80'h10100000010000010010;
mem[2576] = 80'h00109400000208004500;
mem[2577] = 80'h0010002f5fe40000fffd;
mem[2578] = 80'h0010d994c0550102c000;
mem[2579] = 80'h00100001ffabffabffab;
mem[2580] = 80'h0010ff1bb7d64195ad40;
mem[2581] = 80'h001096550cab5d60abda;
mem[2582] = 80'h0010024872b438cb7367;
mem[2583] = 80'h0111ad00000000000000;
mem[2584] = 80'h00000000000000000000;
mem[2585] = 80'h00000000000000000000;
mem[2586] = 80'h00000000000000000000;
mem[2587] = 80'h00000000000000000000;
mem[2588] = 80'h10100000010000010010;
mem[2589] = 80'h00109400000208004500;
mem[2590] = 80'h0010002f5fe50000fffd;
mem[2591] = 80'h0010d993c0550102c000;
mem[2592] = 80'h00100001ffabffabffab;
mem[2593] = 80'h0010ff1ac6086d4dd482;
mem[2594] = 80'h0010299ede2cb0956453;
mem[2595] = 80'h001053f7ea609d6f1566;
mem[2596] = 80'h0111cb00000000000000;
mem[2597] = 80'h10100000010000010010;
mem[2598] = 80'h00109400000208004500;
mem[2599] = 80'h0010002f5fe60000fffd;
mem[2600] = 80'h0010d992c0550102c000;
mem[2601] = 80'h00100001ffabffabffab;
mem[2602] = 80'h0010ff19546a18255ec5;
mem[2603] = 80'h0010e9c2a9a4868b14d8;
mem[2604] = 80'h0010a1b2f7136d6de1ff;
mem[2605] = 80'h01119800000000000000;
mem[2606] = 80'h00000000000000000000;
mem[2607] = 80'h00000000000000000000;
mem[2608] = 80'h00000000000000000000;
mem[2609] = 80'h10100000010000010010;
mem[2610] = 80'h00109400000208004500;
mem[2611] = 80'h0010002f5fe70000fffd;
mem[2612] = 80'h0010d991c0550102c000;
mem[2613] = 80'h00100001ffabffabffab;
mem[2614] = 80'h0010ff1825b434fd2707;
mem[2615] = 80'h001056097b236b7ec4c1;
mem[2616] = 80'h0010f07ad646b6b18d1c;
mem[2617] = 80'h0111e300000000000000;
mem[2618] = 80'h10100000010000010010;
mem[2619] = 80'h00109400000208004500;
mem[2620] = 80'h0010002f5fe80000fffd;
mem[2621] = 80'h0010d990c0550102c000;
mem[2622] = 80'h00100001ffabffabffab;
mem[2623] = 80'h0010ff171de3cd8777da;
mem[2624] = 80'h0010e8b377865ef2d63e;
mem[2625] = 80'h00106aa14d964fbb0d0d;
mem[2626] = 80'h0111be00000000000000;
mem[2627] = 80'h00000000000000000000;
mem[2628] = 80'h00000000000000000000;
mem[2629] = 80'h00000000000000000000;
mem[2630] = 80'h10100000010000010010;
mem[2631] = 80'h00109400000208004500;
mem[2632] = 80'h0010002f5fe90000fffd;
mem[2633] = 80'h0010d98fc0550102c000;
mem[2634] = 80'h00100001ffabffabffab;
mem[2635] = 80'h0010ff166c3de15f0e18;
mem[2636] = 80'h00105778a501b30706b7;
mem[2637] = 80'h00103b71878a2ba1e646;
mem[2638] = 80'h01113b00000000000000;
mem[2639] = 80'h00000000000000000000;
mem[2640] = 80'h10100000010000010010;
mem[2641] = 80'h00109400000208004500;
mem[2642] = 80'h0010002f5fea0000fffd;
mem[2643] = 80'h0010d98ec0550102c000;
mem[2644] = 80'h00100001ffabffabffab;
mem[2645] = 80'h0010ff15fe5f9437845f;
mem[2646] = 80'h00109724d2898519763c;
mem[2647] = 80'h0010c9349aba20f125e4;
mem[2648] = 80'h01119900000000000000;
mem[2649] = 80'h00000000000000000000;
mem[2650] = 80'h00000000000000000000;
mem[2651] = 80'h00000000000000000000;
mem[2652] = 80'h00000000000000000000;
mem[2653] = 80'h10100000010000010010;
mem[2654] = 80'h00109400000208004500;
mem[2655] = 80'h0010002f5feb0000fffd;
mem[2656] = 80'h0010d98dc0550102c000;
mem[2657] = 80'h00100001ffabffabffab;
mem[2658] = 80'h0010ff148f81b8effd9d;
mem[2659] = 80'h001028ef000e68eca645;
mem[2660] = 80'h001098f791b5575d581c;
mem[2661] = 80'h01119700000000000000;
mem[2662] = 80'h00000000000000000000;
mem[2663] = 80'h10100000010000010010;
mem[2664] = 80'h00109400000208004500;
mem[2665] = 80'h0010002f5fec0000fffd;
mem[2666] = 80'h0010d98cc0550102c000;
mem[2667] = 80'h00100001ffabffabffab;
mem[2668] = 80'h0010ff13ab45523ee912;
mem[2669] = 80'h0010a857ef1f04d0477e;
mem[2670] = 80'h00107d6ba12417d9048d;
mem[2671] = 80'h01111800000000000000;
mem[2672] = 80'h00000000000000000000;
mem[2673] = 80'h00000000000000000000;
mem[2674] = 80'h00000000000000000000;
mem[2675] = 80'h10100000010000010010;
mem[2676] = 80'h00109400000208004500;
mem[2677] = 80'h0010002f5fed0000fffd;
mem[2678] = 80'h0010d98bc0550102c000;
mem[2679] = 80'h00100001ffabffabffab;
mem[2680] = 80'h0010ff12da9b7ee690d0;
mem[2681] = 80'h0010179c3d98e9259737;
mem[2682] = 80'h00102cad3f5bd405a26a;
mem[2683] = 80'h01110500000000000000;
mem[2684] = 80'h00000000000000000000;
mem[2685] = 80'h10100000010000010010;
mem[2686] = 80'h00109400000208004500;
mem[2687] = 80'h0010002f5fee0000fffd;
mem[2688] = 80'h0010d98ac0550102c000;
mem[2689] = 80'h00100001ffabffabffab;
mem[2690] = 80'h0010ff1148f90b8e1a97;
mem[2691] = 80'h0010d7c04a10df3be67b;
mem[2692] = 80'h0010de50d1f5f978cdd9;
mem[2693] = 80'h01115f00000000000000;
mem[2694] = 80'h00000000000000000000;
mem[2695] = 80'h10100000010000010010;
mem[2696] = 80'h00109400000208004500;
mem[2697] = 80'h0010002f5fef0000fffd;
mem[2698] = 80'h0010d989c0550102c000;
mem[2699] = 80'h00100001ffabffabffab;
mem[2700] = 80'h0010ff10392727566355;
mem[2701] = 80'h0010680b989732ce363a;
mem[2702] = 80'h00108f1fe6515d2fc6df;
mem[2703] = 80'h01116100000000000000;
mem[2704] = 80'h00000000000000000000;
mem[2705] = 80'h00000000000000000000;
mem[2706] = 80'h00000000000000000000;
mem[2707] = 80'h10100000010000010010;
mem[2708] = 80'h00109400000208004500;
mem[2709] = 80'h0010002f5ff00000fffd;
mem[2710] = 80'h0010d988c0550102c000;
mem[2711] = 80'h00100001ffabffabffab;
mem[2712] = 80'h0010ff0f3856f97abb2c;
mem[2713] = 80'h0010aab4535ab423c396;
mem[2714] = 80'h0010ea92d795db2d1ece;
mem[2715] = 80'h0111f900000000000000;
mem[2716] = 80'h00000000000000000000;
mem[2717] = 80'h10100000010000010010;
mem[2718] = 80'h00109400000208004500;
mem[2719] = 80'h0010002f5ff10000fffd;
mem[2720] = 80'h0010d987c0550102c000;
mem[2721] = 80'h00100001ffabffabffab;
mem[2722] = 80'h0010ff0e4988d5a2c2ee;
mem[2723] = 80'h0010157f81dd59d613d7;
mem[2724] = 80'h0010bbdde0ef7ce8458a;
mem[2725] = 80'h01110900000000000000;
mem[2726] = 80'h00000000000000000000;
mem[2727] = 80'h00000000000000000000;
mem[2728] = 80'h00000000000000000000;
mem[2729] = 80'h10100000010000010010;
mem[2730] = 80'h00109400000208004500;
mem[2731] = 80'h0010002f5ff20000fffd;
mem[2732] = 80'h0010d986c0550102c000;
mem[2733] = 80'h00100001ffabffabffab;
mem[2734] = 80'h0010ff0ddbeaa0ca48a9;
mem[2735] = 80'h0010d523f6556fc86394;
mem[2736] = 80'h0010490700b652b90f97;
mem[2737] = 80'h0111f100000000000000;
mem[2738] = 80'h00000000000000000000;
mem[2739] = 80'h10100000010000010010;
mem[2740] = 80'h00109400000208004500;
mem[2741] = 80'h0010002f5ff30000fffd;
mem[2742] = 80'h0010d985c0550102c000;
mem[2743] = 80'h00100001ffabffabffab;
mem[2744] = 80'h0010ff0caa348c12316b;
mem[2745] = 80'h00106ae824d2823db3d5;
mem[2746] = 80'h00101848372b83e70c7a;
mem[2747] = 80'h0111e100000000000000;
mem[2748] = 80'h00000000000000000000;
mem[2749] = 80'h00000000000000000000;
mem[2750] = 80'h00000000000000000000;
mem[2751] = 80'h00000000000000000000;
mem[2752] = 80'h10100000010000010010;
mem[2753] = 80'h00109400000208004500;
mem[2754] = 80'h0010002f5ff40000fffd;
mem[2755] = 80'h0010d984c0550102c000;
mem[2756] = 80'h00100001ffabffabffab;
mem[2757] = 80'h0010ff0b8ef066c325e4;
mem[2758] = 80'h0010ea50cbc3ee015296;
mem[2759] = 80'h0010fd55f758f99d35ff;
mem[2760] = 80'h0111c300000000000000;
mem[2761] = 80'h10100000010000010010;
mem[2762] = 80'h00109400000208004500;
mem[2763] = 80'h0010002f5ff50000fffd;
mem[2764] = 80'h0010d983c0550102c000;
mem[2765] = 80'h00100001ffabffabffab;
mem[2766] = 80'h0010ff0aff2e4a1b5c26;
mem[2767] = 80'h0010559b194403f48296;
mem[2768] = 80'h0010ac243df67bf2bda7;
mem[2769] = 80'h01118400000000000000;
mem[2770] = 80'h00000000000000000000;
mem[2771] = 80'h00000000000000000000;
mem[2772] = 80'h00000000000000000000;
mem[2773] = 80'h10100000010000010010;
mem[2774] = 80'h00109400000208004500;
mem[2775] = 80'h0010002f5ff60000fffd;
mem[2776] = 80'h0010d982c0550102c000;
mem[2777] = 80'h00100001ffabffabffab;
mem[2778] = 80'h0010ff096d4c3f73d661;
mem[2779] = 80'h001095c76ecc35eaf215;
mem[2780] = 80'h00105ee8895868535c00;
mem[2781] = 80'h01117000000000000000;
mem[2782] = 80'h00000000000000000000;
mem[2783] = 80'h10100000010000010010;
mem[2784] = 80'h00109400000208004500;
mem[2785] = 80'h0010002f5ff70000fffd;
mem[2786] = 80'h0010d981c0550102c000;
mem[2787] = 80'h00100001ffabffabffab;
mem[2788] = 80'h0010ff081c9213abafa3;
mem[2789] = 80'h00102a0cbc4bd81f2194;
mem[2790] = 80'h00100fe8ba2276990177;
mem[2791] = 80'h01119e00000000000000;
mem[2792] = 80'h00000000000000000000;
mem[2793] = 80'h00000000000000000000;
mem[2794] = 80'h00000000000000000000;
mem[2795] = 80'h10100000010000010010;
mem[2796] = 80'h00109400000208004500;
mem[2797] = 80'h0010002f5ff80000fffd;
mem[2798] = 80'h0010d980c0550102c000;
mem[2799] = 80'h00100001ffabffabffab;
mem[2800] = 80'h0010ff0724c5ead1ff7e;
mem[2801] = 80'h001094b6b0eeed933372;
mem[2802] = 80'h0010958acaac2a2ccbf6;
mem[2803] = 80'h0111a000000000000000;
mem[2804] = 80'h00000000000000000000;
mem[2805] = 80'h10100000010000010010;
mem[2806] = 80'h00109400000208004500;
mem[2807] = 80'h0010002f5ff90000fffd;
mem[2808] = 80'h0010d97fc0550102c000;
mem[2809] = 80'h00100001ffabffabffab;
mem[2810] = 80'h0010ff06551bc60986bc;
mem[2811] = 80'h00102b7d62690066e373;
mem[2812] = 80'h0010c4c8318ef6277c1a;
mem[2813] = 80'h01112c00000000000000;
mem[2814] = 80'h00000000000000000000;
mem[2815] = 80'h00000000000000000000;
mem[2816] = 80'h00000000000000000000;
mem[2817] = 80'h00000000000000000000;
mem[2818] = 80'h10100000010000010010;
mem[2819] = 80'h00109400000208004500;
mem[2820] = 80'h0010002f5ffa0000fffd;
mem[2821] = 80'h0010d97ec0550102c000;
mem[2822] = 80'h00100001ffabffabffab;
mem[2823] = 80'h0010ff05c779b3610cfb;
mem[2824] = 80'h0010eb2115e1367893f0;
mem[2825] = 80'h0010360485b3f122900b;
mem[2826] = 80'h01119800000000000000;
mem[2827] = 80'h10100000010000010010;
mem[2828] = 80'h00109400000208004500;
mem[2829] = 80'h0010002f5ffb0000fffd;
mem[2830] = 80'h0010d97dc0550102c000;
mem[2831] = 80'h00100001ffabffabffab;
mem[2832] = 80'h0010ff04b6a79fb97539;
mem[2833] = 80'h001054eac766db8d4372;
mem[2834] = 80'h00106708b506dd3b3e25;
mem[2835] = 80'h01110d00000000000000;
mem[2836] = 80'h00000000000000000000;
mem[2837] = 80'h00000000000000000000;
mem[2838] = 80'h00000000000000000000;
mem[2839] = 80'h10100000010000010010;
mem[2840] = 80'h00109400000208004500;
mem[2841] = 80'h0010002f5ffc0000fffd;
mem[2842] = 80'h0010d97cc0550102c000;
mem[2843] = 80'h00100001ffabffabffab;
mem[2844] = 80'h0010ff039263756861b6;
mem[2845] = 80'h0010d4522877b7b1a231;
mem[2846] = 80'h0010821575b748644dd9;
mem[2847] = 80'h0111e600000000000000;
mem[2848] = 80'h00000000000000000000;
mem[2849] = 80'h10100000010000010010;
mem[2850] = 80'h00109400000208004500;
mem[2851] = 80'h0010002f5ffd0000fffd;
mem[2852] = 80'h0010d97bc0550102c000;
mem[2853] = 80'h00100001ffabffabffab;
mem[2854] = 80'h0010ff02e3bd59b01874;
mem[2855] = 80'h00106b99faf05a447270;
mem[2856] = 80'h0010d35a428161a109f1;
mem[2857] = 80'h01113000000000000000;
mem[2858] = 80'h00000000000000000000;
mem[2859] = 80'h00000000000000000000;
mem[2860] = 80'h00000000000000000000;
mem[2861] = 80'h10100000010000010010;
mem[2862] = 80'h00109400000208004500;
mem[2863] = 80'h0010002f5ffe0000fffd;
mem[2864] = 80'h0010d97ac0550102c000;
mem[2865] = 80'h00100001ffabffabffab;
mem[2866] = 80'h0010ff0171df2cd89233;
mem[2867] = 80'h0010abc58d786c5a02b3;
mem[2868] = 80'h0010219b3a2ccb7e0d41;
mem[2869] = 80'h01113800000000000000;
mem[2870] = 80'h00000000000000000000;
mem[2871] = 80'h00000000000000000000;
mem[2872] = 80'h00000000000000000000;
mem[2873] = 80'h10100000010000010010;
mem[2874] = 80'h00109400000208004500;
mem[2875] = 80'h0010002f5fff0000fffd;
mem[2876] = 80'h0010d979c0550102c000;
mem[2877] = 80'h00100001ffabffabffab;
mem[2878] = 80'h0010ff0000010000ebf1;
mem[2879] = 80'h0010140e5fff81afd2f2;
mem[2880] = 80'h001070d40d88cdedc49f;
mem[2881] = 80'h01113e00000000000000;
mem[2882] = 80'h00000000000000000000;
mem[2883] = 80'h10100000010000010010;
mem[2884] = 80'h00109400000208004500;
mem[2885] = 80'h0010002f60000000fffd;
mem[2886] = 80'h0010d978c0550102c000;
mem[2887] = 80'h00100001ffabffabffab;
mem[2888] = 80'h0010ffff2f4b1bb73cb0;
mem[2889] = 80'h00108148d182dafc9cd2;
mem[2890] = 80'h0010bf7d873566a9f166;
mem[2891] = 80'h0111e200000000000000;
mem[2892] = 80'h00000000000000000000;
mem[2893] = 80'h00000000000000000000;
mem[2894] = 80'h00000000000000000000;
mem[2895] = 80'h10100000010000010010;
mem[2896] = 80'h00109400000208004500;
mem[2897] = 80'h0010002f60010000fffd;
mem[2898] = 80'h0010d977c0550102c000;
mem[2899] = 80'h00100001ffabffabffab;
mem[2900] = 80'h0010fffe5e95376f4572;
mem[2901] = 80'h00103e83030537094c92;
mem[2902] = 80'h0010ee018164ef8751ef;
mem[2903] = 80'h0111b400000000000000;
mem[2904] = 80'h00000000000000000000;
mem[2905] = 80'h10100000010000010010;
mem[2906] = 80'h00109400000208004500;
mem[2907] = 80'h0010002f60020000fffd;
mem[2908] = 80'h0010d976c0550102c000;
mem[2909] = 80'h00100001ffabffabffab;
mem[2910] = 80'h0010fffdccf74207cf35;
mem[2911] = 80'h0010fedf748d01173c51;
mem[2912] = 80'h00101cc0f9375a9e9468;
mem[2913] = 80'h0111bb00000000000000;
mem[2914] = 80'h00000000000000000000;
mem[2915] = 80'h00000000000000000000;
mem[2916] = 80'h00000000000000000000;
mem[2917] = 80'h10100000010000010010;
mem[2918] = 80'h00109400000208004500;
mem[2919] = 80'h0010002f60030000fffd;
mem[2920] = 80'h0010d975c0550102c000;
mem[2921] = 80'h00100001ffabffabffab;
mem[2922] = 80'h0010fffcbd296edfb6f7;
mem[2923] = 80'h00104114a60aece2ec10;
mem[2924] = 80'h00104d8fce60403cb326;
mem[2925] = 80'h01119600000000000000;
mem[2926] = 80'h00000000000000000000;
mem[2927] = 80'h10100000010000010010;
mem[2928] = 80'h00109400000208004500;
mem[2929] = 80'h0010002f60040000fffd;
mem[2930] = 80'h0010d974c0550102c000;
mem[2931] = 80'h00100001ffabffabffab;
mem[2932] = 80'h0010fffb99ed840ea278;
mem[2933] = 80'h0010c1ac491b80de0d53;
mem[2934] = 80'h0010a8920e03ef4cbed8;
mem[2935] = 80'h01110800000000000000;
mem[2936] = 80'h00000000000000000000;
mem[2937] = 80'h00000000000000000000;
mem[2938] = 80'h00000000000000000000;
mem[2939] = 80'h00000000000000000000;
mem[2940] = 80'h10100000010000010010;
mem[2941] = 80'h00109400000208004500;
mem[2942] = 80'h0010002f60050000fffd;
mem[2943] = 80'h0010d973c0550102c000;
mem[2944] = 80'h00100001ffabffabffab;
mem[2945] = 80'h0010fffae833a8d6dbba;
mem[2946] = 80'h00107e679b9c6d2bddd2;
mem[2947] = 80'h0010f9cb6d71c613e0ca;
mem[2948] = 80'h01114500000000000000;
mem[2949] = 80'h10100000010000010010;
mem[2950] = 80'h00109400000208004500;
mem[2951] = 80'h0010002f60060000fffd;
mem[2952] = 80'h0010d972c0550102c000;
mem[2953] = 80'h00100001ffabffabffab;
mem[2954] = 80'h0010fff97a51ddbe51fd;
mem[2955] = 80'h0010be3bec145b35ad51;
mem[2956] = 80'h00100b07d919beaac9ad;
mem[2957] = 80'h0111f600000000000000;
mem[2958] = 80'h00000000000000000000;
mem[2959] = 80'h00000000000000000000;
mem[2960] = 80'h00000000000000000000;
mem[2961] = 80'h10100000010000010010;
mem[2962] = 80'h00109400000208004500;
mem[2963] = 80'h0010002f60070000fffd;
mem[2964] = 80'h0010d971c0550102c000;
mem[2965] = 80'h00100001ffabffabffab;
mem[2966] = 80'h0010fff80b8ff166283f;
mem[2967] = 80'h001001f03e93b6c07d57;
mem[2968] = 80'h00105adcb55a55a17661;
mem[2969] = 80'h01117f00000000000000;
mem[2970] = 80'h10100000010000010010;
mem[2971] = 80'h00109400000208004500;
mem[2972] = 80'h0010002f60080000fffd;
mem[2973] = 80'h0010d970c0550102c000;
mem[2974] = 80'h00100001ffabffabffab;
mem[2975] = 80'h0010fff733d8081c78e2;
mem[2976] = 80'h0010bf4a3236834c6fa9;
mem[2977] = 80'h0010c0341f86863c7b15;
mem[2978] = 80'h01115900000000000000;
mem[2979] = 80'h00000000000000000000;
mem[2980] = 80'h00000000000000000000;
mem[2981] = 80'h00000000000000000000;
mem[2982] = 80'h10100000010000010010;
mem[2983] = 80'h00109400000208004500;
mem[2984] = 80'h0010002f60090000fffd;
mem[2985] = 80'h0010d96fc0550102c000;
mem[2986] = 80'h00100001ffabffabffab;
mem[2987] = 80'h0010fff6420624c40120;
mem[2988] = 80'h00100081e0b16eb9b830;
mem[2989] = 80'h00109162369fc72f0bca;
mem[2990] = 80'h01114f00000000000000;
mem[2991] = 80'h00000000000000000000;
mem[2992] = 80'h10100000010000010010;
mem[2993] = 80'h00109400000208004500;
mem[2994] = 80'h0010002f600a0000fffd;
mem[2995] = 80'h0010d96ec0550102c000;
mem[2996] = 80'h00100001ffabffabffab;
mem[2997] = 80'h0010fff5d06451ac8b67;
mem[2998] = 80'h0010c0dd973958a7c8bb;
mem[2999] = 80'h001063272bf0494bfe99;
mem[3000] = 80'h01114d00000000000000;
mem[3001] = 80'h00000000000000000000;
mem[3002] = 80'h00000000000000000000;
mem[3003] = 80'h00000000000000000000;
mem[3004] = 80'h00000000000000000000;
mem[3005] = 80'h10100000010000010010;
mem[3006] = 80'h00109400000208004500;
mem[3007] = 80'h0010002f600b0000fffd;
mem[3008] = 80'h0010d96dc0550102c000;
mem[3009] = 80'h00100001ffabffabffab;
mem[3010] = 80'h0010fff4a1ba7d74f2a5;
mem[3011] = 80'h00107f1645beb55218b2;
mem[3012] = 80'h001032ec7970ae36a48e;
mem[3013] = 80'h0111a200000000000000;
mem[3014] = 80'h00000000000000000000;
mem[3015] = 80'h10100000010000010010;
mem[3016] = 80'h00109400000208004500;
mem[3017] = 80'h0010002f600c0000fffd;
mem[3018] = 80'h0010d96cc0550102c000;
mem[3019] = 80'h00100001ffabffabffab;
mem[3020] = 80'h0010fff3857e97a5e62a;
mem[3021] = 80'h0010ffaeaaafd96ef9c9;
mem[3022] = 80'h0010d77d85a8214a6ef8;
mem[3023] = 80'h01116200000000000000;
mem[3024] = 80'h00000000000000000000;
mem[3025] = 80'h00000000000000000000;
mem[3026] = 80'h00000000000000000000;
mem[3027] = 80'h10100000010000010010;
mem[3028] = 80'h00109400000208004500;
mem[3029] = 80'h0010002f600d0000fffd;
mem[3030] = 80'h0010d96bc0550102c000;
mem[3031] = 80'h00100001ffabffabffab;
mem[3032] = 80'h0010fff2f4a0bb7d9fe8;
mem[3033] = 80'h001040657828349b29b0;
mem[3034] = 80'h001086be8e6e832d01d1;
mem[3035] = 80'h0111b800000000000000;
mem[3036] = 80'h00000000000000000000;
mem[3037] = 80'h10100000010000010010;
mem[3038] = 80'h00109400000208004500;
mem[3039] = 80'h0010002f600e0000fffd;
mem[3040] = 80'h0010d96ac0550102c000;
mem[3041] = 80'h00100001ffabffabffab;
mem[3042] = 80'h0010fff166c2ce1515af;
mem[3043] = 80'h001080390fa0028559fa;
mem[3044] = 80'h001074def64f5de05c57;
mem[3045] = 80'h0111bc00000000000000;
mem[3046] = 80'h00000000000000000000;
mem[3047] = 80'h10100000010000010010;
mem[3048] = 80'h00109400000208004500;
mem[3049] = 80'h0010002f600f0000fffd;
mem[3050] = 80'h0010d969c0550102c000;
mem[3051] = 80'h00100001ffabffabffab;
mem[3052] = 80'h0010fff0171ce2cd6c6d;
mem[3053] = 80'h00103ff2dd27ef7089b3;
mem[3054] = 80'h001025186861754ef598;
mem[3055] = 80'h01110d00000000000000;
mem[3056] = 80'h00000000000000000000;
mem[3057] = 80'h00000000000000000000;
mem[3058] = 80'h00000000000000000000;
mem[3059] = 80'h10100000010000010010;
mem[3060] = 80'h00109400000208004500;
mem[3061] = 80'h0010002f60100000fffd;
mem[3062] = 80'h0010d968c0550102c000;
mem[3063] = 80'h00100001ffabffabffab;
mem[3064] = 80'h0010ffef166d3ce1b414;
mem[3065] = 80'h0010fd4d16ea699d7c07;
mem[3066] = 80'h0010401f83b13a42e6e0;
mem[3067] = 80'h0111b400000000000000;
mem[3068] = 80'h00000000000000000000;
mem[3069] = 80'h10100000010000010010;
mem[3070] = 80'h00109400000208004500;
mem[3071] = 80'h0010002f60110000fffd;
mem[3072] = 80'h0010d967c0550102c000;
mem[3073] = 80'h00100001ffabffabffab;
mem[3074] = 80'h0010ffee67b31039cdd6;
mem[3075] = 80'h00104286c46d8468ac5e;
mem[3076] = 80'h001011da6eb901d31f6b;
mem[3077] = 80'h01114d00000000000000;
mem[3078] = 80'h00000000000000000000;
mem[3079] = 80'h00000000000000000000;
mem[3080] = 80'h00000000000000000000;
mem[3081] = 80'h10100000010000010010;
mem[3082] = 80'h00109400000208004500;
mem[3083] = 80'h0010002f60120000fffd;
mem[3084] = 80'h0010d966c0550102c000;
mem[3085] = 80'h00100001ffabffabffab;
mem[3086] = 80'h0010ffedf5d165514791;
mem[3087] = 80'h001082dab3e5b276dd15;
mem[3088] = 80'h0010e3be17529b22ddc2;
mem[3089] = 80'h0111ea00000000000000;
mem[3090] = 80'h00000000000000000000;
mem[3091] = 80'h10100000010000010010;
mem[3092] = 80'h00109400000208004500;
mem[3093] = 80'h0010002f60130000fffd;
mem[3094] = 80'h0010d965c0550102c000;
mem[3095] = 80'h00100001ffabffabffab;
mem[3096] = 80'h0010ffec840f49893e53;
mem[3097] = 80'h00103d1161625f830d5c;
mem[3098] = 80'h0010b278895bac1ccbc0;
mem[3099] = 80'h01110c00000000000000;
mem[3100] = 80'h00000000000000000000;
mem[3101] = 80'h00000000000000000000;
mem[3102] = 80'h00000000000000000000;
mem[3103] = 80'h00000000000000000000;
mem[3104] = 80'h10100000010000010010;
mem[3105] = 80'h00109400000208004500;
mem[3106] = 80'h0010002f60140000fffd;
mem[3107] = 80'h0010d964c0550102c000;
mem[3108] = 80'h00100001ffabffabffab;
mem[3109] = 80'h0010ffeba0cba3582adc;
mem[3110] = 80'h0010bda98e7333bfec64;
mem[3111] = 80'h001057b1ea20e22ebcc5;
mem[3112] = 80'h0111d400000000000000;
mem[3113] = 80'h10100000010000010010;
mem[3114] = 80'h00109400000208004500;
mem[3115] = 80'h0010002f60150000fffd;
mem[3116] = 80'h0010d963c0550102c000;
mem[3117] = 80'h00100001ffabffabffab;
mem[3118] = 80'h0010ffead1158f80531e;
mem[3119] = 80'h001002625cf4de4a3c1d;
mem[3120] = 80'h00100672e12feab8f5d7;
mem[3121] = 80'h01112200000000000000;
mem[3122] = 80'h00000000000000000000;
mem[3123] = 80'h00000000000000000000;
mem[3124] = 80'h00000000000000000000;
mem[3125] = 80'h10100000010000010010;
mem[3126] = 80'h00109400000208004500;
mem[3127] = 80'h0010002f60160000fffd;
mem[3128] = 80'h0010d962c0550102c000;
mem[3129] = 80'h00100001ffabffabffab;
mem[3130] = 80'h0010ffe94377fae8d959;
mem[3131] = 80'h0010c23e2b7ce8544c96;
mem[3132] = 80'h0010f437fc7dd4eefb0d;
mem[3133] = 80'h01118100000000000000;
mem[3134] = 80'h00000000000000000000;
mem[3135] = 80'h10100000010000010010;
mem[3136] = 80'h00109400000208004500;
mem[3137] = 80'h0010002f60170000fffd;
mem[3138] = 80'h0010d961c0550102c000;
mem[3139] = 80'h00100001ffabffabffab;
mem[3140] = 80'h0010ffe832a9d630a09b;
mem[3141] = 80'h00107df5f9fb05a19c1f;
mem[3142] = 80'h0010a5e73608602b991b;
mem[3143] = 80'h01119f00000000000000;
mem[3144] = 80'h00000000000000000000;
mem[3145] = 80'h00000000000000000000;
mem[3146] = 80'h00000000000000000000;
mem[3147] = 80'h10100000010000010010;
mem[3148] = 80'h00109400000208004500;
mem[3149] = 80'h0010002f60180000fffd;
mem[3150] = 80'h0010d960c0550102c000;
mem[3151] = 80'h00100001ffabffabffab;
mem[3152] = 80'h0010ffe70afe2f4af046;
mem[3153] = 80'h0010c34ff55e302d8ee1;
mem[3154] = 80'h00103f0f9cbc8199249c;
mem[3155] = 80'h0111dc00000000000000;
mem[3156] = 80'h00000000000000000000;
mem[3157] = 80'h10100000010000010010;
mem[3158] = 80'h00109400000208004500;
mem[3159] = 80'h0010002f60190000fffd;
mem[3160] = 80'h0010d95fc0550102c000;
mem[3161] = 80'h00100001ffabffabffab;
mem[3162] = 80'h0010ffe67b2003928984;
mem[3163] = 80'h00107c8427d9ddd85ef8;
mem[3164] = 80'h00106ec7bdebe9ed8163;
mem[3165] = 80'h01117700000000000000;
mem[3166] = 80'h00000000000000000000;
mem[3167] = 80'h00000000000000000000;
mem[3168] = 80'h00000000000000000000;
mem[3169] = 80'h00000000000000000000;
mem[3170] = 80'h10100000010000010010;
mem[3171] = 80'h00109400000208004500;
mem[3172] = 80'h0010002f601a0000fffd;
mem[3173] = 80'h0010d95ec0550102c000;
mem[3174] = 80'h00100001ffabffabffab;
mem[3175] = 80'h0010ffe5e94276fa03c3;
mem[3176] = 80'h0010bcd85051ebc62e72;
mem[3177] = 80'h00109cb191054690c6aa;
mem[3178] = 80'h01111700000000000000;
mem[3179] = 80'h10100000010000010010;
mem[3180] = 80'h00109400000208004500;
mem[3181] = 80'h0010002f601b0000fffd;
mem[3182] = 80'h0010d95dc0550102c000;
mem[3183] = 80'h00100001ffabffabffab;
mem[3184] = 80'h0010ffe4989c5a227a01;
mem[3185] = 80'h0010031382d60633fdfb;
mem[3186] = 80'h0010cd380b0a30b0e257;
mem[3187] = 80'h01114200000000000000;
mem[3188] = 80'h00000000000000000000;
mem[3189] = 80'h00000000000000000000;
mem[3190] = 80'h00000000000000000000;
mem[3191] = 80'h10100000010000010010;
mem[3192] = 80'h00109400000208004500;
mem[3193] = 80'h0010002f601c0000fffd;
mem[3194] = 80'h0010d95cc0550102c000;
mem[3195] = 80'h00100001ffabffabffab;
mem[3196] = 80'h0010ffe3bc58b0f36e8e;
mem[3197] = 80'h001083ab6dc76a0f1c80;
mem[3198] = 80'h001028a9f7958bbb05ad;
mem[3199] = 80'h01111c00000000000000;
mem[3200] = 80'h00000000000000000000;
mem[3201] = 80'h10100000010000010010;
mem[3202] = 80'h00109400000208004500;
mem[3203] = 80'h0010002f601d0000fffd;
mem[3204] = 80'h0010d95bc0550102c000;
mem[3205] = 80'h00100001ffabffabffab;
mem[3206] = 80'h0010ffe2cd869c2b174c;
mem[3207] = 80'h00103c60bf4087faccf9;
mem[3208] = 80'h0010796afc1eb846f85b;
mem[3209] = 80'h01110400000000000000;
mem[3210] = 80'h00000000000000000000;
mem[3211] = 80'h00000000000000000000;
mem[3212] = 80'h00000000000000000000;
mem[3213] = 80'h10100000010000010010;
mem[3214] = 80'h00109400000208004500;
mem[3215] = 80'h0010002f601e0000fffd;
mem[3216] = 80'h0010d95ac0550102c000;
mem[3217] = 80'h00100001ffabffabffab;
mem[3218] = 80'h0010ffe15fe4e9439d0b;
mem[3219] = 80'h0010fc3cc8c8b1e4bc32;
mem[3220] = 80'h00108b222dab2dce543d;
mem[3221] = 80'h01119200000000000000;
mem[3222] = 80'h00000000000000000000;
mem[3223] = 80'h00000000000000000000;
mem[3224] = 80'h00000000000000000000;
mem[3225] = 80'h10100000010000010010;
mem[3226] = 80'h00109400000208004500;
mem[3227] = 80'h0010002f601f0000fffd;
mem[3228] = 80'h0010d959c0550102c000;
mem[3229] = 80'h00100001ffabffabffab;
mem[3230] = 80'h0010ffe02e3ac59be4c9;
mem[3231] = 80'h001043f71a4f5c116c7b;
mem[3232] = 80'h0010dae4b3c771c265d5;
mem[3233] = 80'h0111b600000000000000;
mem[3234] = 80'h00000000000000000000;
mem[3235] = 80'h10100000010000010010;
mem[3236] = 80'h00109400000208004500;
mem[3237] = 80'h0010002f60200000fffd;
mem[3238] = 80'h0010d958c0550102c000;
mem[3239] = 80'h00100001ffabffabffab;
mem[3240] = 80'h0010ffdf5d07551a2df8;
mem[3241] = 80'h001079435f53bc3f575d;
mem[3242] = 80'h001041b46c1e853ac4fa;
mem[3243] = 80'h0111f400000000000000;
mem[3244] = 80'h00000000000000000000;
mem[3245] = 80'h00000000000000000000;
mem[3246] = 80'h00000000000000000000;
mem[3247] = 80'h10100000010000010010;
mem[3248] = 80'h00109400000208004500;
mem[3249] = 80'h0010002f60210000fffd;
mem[3250] = 80'h0010d957c0550102c000;
mem[3251] = 80'h00100001ffabffabffab;
mem[3252] = 80'h0010ffde2cd979c2543a;
mem[3253] = 80'h0010c6888dd451ca871c;
mem[3254] = 80'h001010fb5b0c6b64879a;
mem[3255] = 80'h0111a600000000000000;
mem[3256] = 80'h00000000000000000000;
mem[3257] = 80'h10100000010000010010;
mem[3258] = 80'h00109400000208004500;
mem[3259] = 80'h0010002f60220000fffd;
mem[3260] = 80'h0010d956c0550102c000;
mem[3261] = 80'h00100001ffabffabffab;
mem[3262] = 80'h0010ffddbebb0caade7d;
mem[3263] = 80'h001006d4fa5c67d4f7cf;
mem[3264] = 80'h0010e239502fc2b81cf7;
mem[3265] = 80'h0111d500000000000000;
mem[3266] = 80'h00000000000000000000;
mem[3267] = 80'h00000000000000000000;
mem[3268] = 80'h00000000000000000000;
mem[3269] = 80'h10100000010000010010;
mem[3270] = 80'h00109400000208004500;
mem[3271] = 80'h0010002f60230000fffd;
mem[3272] = 80'h0010d955c0550102c000;
mem[3273] = 80'h00100001ffabffabffab;
mem[3274] = 80'h0010ffdccf652072a7bf;
mem[3275] = 80'h0010b91f28db8a21278e;
mem[3276] = 80'h0010b376676ab9071af8;
mem[3277] = 80'h0111ba00000000000000;
mem[3278] = 80'h00000000000000000000;
mem[3279] = 80'h10100000010000010010;
mem[3280] = 80'h00109400000208004500;
mem[3281] = 80'h0010002f60240000fffd;
mem[3282] = 80'h0010d954c0550102c000;
mem[3283] = 80'h00100001ffabffabffab;
mem[3284] = 80'h0010ffdbeba1caa3b330;
mem[3285] = 80'h001039a7c7cae61dc73d;
mem[3286] = 80'h0010564f56913aa548f5;
mem[3287] = 80'h01118700000000000000;
mem[3288] = 80'h00000000000000000000;
mem[3289] = 80'h00000000000000000000;
mem[3290] = 80'h00000000000000000000;
mem[3291] = 80'h00000000000000000000;
mem[3292] = 80'h10100000010000010010;
mem[3293] = 80'h00109400000208004500;
mem[3294] = 80'h0010002f60250000fffd;
mem[3295] = 80'h0010d953c0550102c000;
mem[3296] = 80'h00100001ffabffabffab;
mem[3297] = 80'h0010ffda9a7fe67bcaf2;
mem[3298] = 80'h0010866c154d0be8177c;
mem[3299] = 80'h0010070061198c83012b;
mem[3300] = 80'h01114b00000000000000;
mem[3301] = 80'h10100000010000010010;
mem[3302] = 80'h00109400000208004500;
mem[3303] = 80'h0010002f60260000fffd;
mem[3304] = 80'h0010d952c0550102c000;
mem[3305] = 80'h00100001ffabffabffab;
mem[3306] = 80'h0010ffd9081d931340b5;
mem[3307] = 80'h0010463062c53df667cf;
mem[3308] = 80'h0010f5c940bb9e3c1242;
mem[3309] = 80'h0111ac00000000000000;
mem[3310] = 80'h00000000000000000000;
mem[3311] = 80'h00000000000000000000;
mem[3312] = 80'h00000000000000000000;
mem[3313] = 80'h10100000010000010010;
mem[3314] = 80'h00109400000208004500;
mem[3315] = 80'h0010002f60270000fffd;
mem[3316] = 80'h0010d951c0550102c000;
mem[3317] = 80'h00100001ffabffabffab;
mem[3318] = 80'h0010ffd879c3bfcb3977;
mem[3319] = 80'h0010f9fbb042d003b7cf;
mem[3320] = 80'h0010a4b88a562b0d7ba3;
mem[3321] = 80'h0111b000000000000000;
mem[3322] = 80'h10100000010000010010;
mem[3323] = 80'h00109400000208004500;
mem[3324] = 80'h0010002f60280000fffd;
mem[3325] = 80'h0010d950c0550102c000;
mem[3326] = 80'h00100001ffabffabffab;
mem[3327] = 80'h0010ffd7419446b169aa;
mem[3328] = 80'h00104741bce7e58fa539;
mem[3329] = 80'h00103ed9896cb65e533c;
mem[3330] = 80'h0111a500000000000000;
mem[3331] = 80'h00000000000000000000;
mem[3332] = 80'h00000000000000000000;
mem[3333] = 80'h00000000000000000000;
mem[3334] = 80'h10100000010000010010;
mem[3335] = 80'h00109400000208004500;
mem[3336] = 80'h0010002f60290000fffd;
mem[3337] = 80'h0010d94fc0550102c000;
mem[3338] = 80'h00100001ffabffabffab;
mem[3339] = 80'h0010ffd6304a6a691068;
mem[3340] = 80'h0010f88a6e60087a75b8;
mem[3341] = 80'h00106f80ea6f15fafc86;
mem[3342] = 80'h01114200000000000000;
mem[3343] = 80'h00000000000000000000;
mem[3344] = 80'h10100000010000010010;
mem[3345] = 80'h00109400000208004500;
mem[3346] = 80'h0010002f602a0000fffd;
mem[3347] = 80'h0010d94ec0550102c000;
mem[3348] = 80'h00100001ffabffabffab;
mem[3349] = 80'h0010ffd5a2281f019a2f;
mem[3350] = 80'h001038d619e83e64052b;
mem[3351] = 80'h00109d4f2d3443c0c688;
mem[3352] = 80'h01119e00000000000000;
mem[3353] = 80'h00000000000000000000;
mem[3354] = 80'h00000000000000000000;
mem[3355] = 80'h00000000000000000000;
mem[3356] = 80'h00000000000000000000;
mem[3357] = 80'h10100000010000010010;
mem[3358] = 80'h00109400000208004500;
mem[3359] = 80'h0010002f602b0000fffd;
mem[3360] = 80'h0010d94dc0550102c000;
mem[3361] = 80'h00100001ffabffabffab;
mem[3362] = 80'h0010ffd4d3f633d9e3ed;
mem[3363] = 80'h0010871dcb6fd391d52a;
mem[3364] = 80'h0010cc0dd61576debff5;
mem[3365] = 80'h01110400000000000000;
mem[3366] = 80'h00000000000000000000;
mem[3367] = 80'h10100000010000010010;
mem[3368] = 80'h00109400000208004500;
mem[3369] = 80'h0010002f602c0000fffd;
mem[3370] = 80'h0010d94cc0550102c000;
mem[3371] = 80'h00100001ffabffabffab;
mem[3372] = 80'h0010ffd3f732d908f762;
mem[3373] = 80'h001007a5247ebfad3459;
mem[3374] = 80'h00102915834e6b715187;
mem[3375] = 80'h01116000000000000000;
mem[3376] = 80'h00000000000000000000;
mem[3377] = 80'h00000000000000000000;
mem[3378] = 80'h00000000000000000000;
mem[3379] = 80'h10100000010000010010;
mem[3380] = 80'h00109400000208004500;
mem[3381] = 80'h0010002f602d0000fffd;
mem[3382] = 80'h0010d94bc0550102c000;
mem[3383] = 80'h00100001ffabffabffab;
mem[3384] = 80'h0010ffd286ecf5d08ea0;
mem[3385] = 80'h0010b86ef6f95258ebdb;
mem[3386] = 80'h0010783582fd0b0ae2cc;
mem[3387] = 80'h0111dd00000000000000;
mem[3388] = 80'h00000000000000000000;
mem[3389] = 80'h10100000010000010010;
mem[3390] = 80'h00109400000208004500;
mem[3391] = 80'h0010002f602e0000fffd;
mem[3392] = 80'h0010d94ac0550102c000;
mem[3393] = 80'h00100001ffabffabffab;
mem[3394] = 80'h0010ffd1148e80b804e7;
mem[3395] = 80'h00107832817164469b68;
mem[3396] = 80'h00108afca3b13d06cb5b;
mem[3397] = 80'h0111c600000000000000;
mem[3398] = 80'h00000000000000000000;
mem[3399] = 80'h10100000010000010010;
mem[3400] = 80'h00109400000208004500;
mem[3401] = 80'h0010002f602f0000fffd;
mem[3402] = 80'h0010d949c0550102c000;
mem[3403] = 80'h00100001ffabffabffab;
mem[3404] = 80'h0010ffd06550ac607d25;
mem[3405] = 80'h0010c7f953f689b34b29;
mem[3406] = 80'h0010dbb394d80f235f65;
mem[3407] = 80'h01119f00000000000000;
mem[3408] = 80'h00000000000000000000;
mem[3409] = 80'h00000000000000000000;
mem[3410] = 80'h00000000000000000000;
mem[3411] = 80'h10100000010000010010;
mem[3412] = 80'h00109400000208004500;
mem[3413] = 80'h0010002f60300000fffd;
mem[3414] = 80'h0010d948c0550102c000;
mem[3415] = 80'h00100001ffabffabffab;
mem[3416] = 80'h0010ffcf6421724ca55c;
mem[3417] = 80'h00100546983b0f5ebe95;
mem[3418] = 80'h0010be3dd6b2832484f1;
mem[3419] = 80'h01119000000000000000;
mem[3420] = 80'h00000000000000000000;
mem[3421] = 80'h10100000010000010010;
mem[3422] = 80'h00109400000208004500;
mem[3423] = 80'h0010002f60310000fffd;
mem[3424] = 80'h0010d947c0550102c000;
mem[3425] = 80'h00100001ffabffabffab;
mem[3426] = 80'h0010ffce15ff5e94dc9e;
mem[3427] = 80'h0010ba8d4abce2ab6ed4;
mem[3428] = 80'h0010ef72e1c1866ca6af;
mem[3429] = 80'h01118900000000000000;
mem[3430] = 80'h00000000000000000000;
mem[3431] = 80'h00000000000000000000;
mem[3432] = 80'h00000000000000000000;
mem[3433] = 80'h10100000010000010010;
mem[3434] = 80'h00109400000208004500;
mem[3435] = 80'h0010002f60320000fffd;
mem[3436] = 80'h0010d946c0550102c000;
mem[3437] = 80'h00100001ffabffabffab;
mem[3438] = 80'h0010ffcd879d2bfc56d9;
mem[3439] = 80'h00107ad13d34d4b51e87;
mem[3440] = 80'h00101dab72d1b9ff436d;
mem[3441] = 80'h01117d00000000000000;
mem[3442] = 80'h00000000000000000000;
mem[3443] = 80'h10100000010000010010;
mem[3444] = 80'h00109400000208004500;
mem[3445] = 80'h0010002f60330000fffd;
mem[3446] = 80'h0010d945c0550102c000;
mem[3447] = 80'h00100001ffabffabffab;
mem[3448] = 80'h0010ffccf64307242f1b;
mem[3449] = 80'h0010c51aefb33940cec7;
mem[3450] = 80'h00104cd7740255766579;
mem[3451] = 80'h01115700000000000000;
mem[3452] = 80'h00000000000000000000;
mem[3453] = 80'h00000000000000000000;
mem[3454] = 80'h00000000000000000000;
mem[3455] = 80'h00000000000000000000;
mem[3456] = 80'h10100000010000010010;
mem[3457] = 80'h00109400000208004500;
mem[3458] = 80'h0010002f60340000fffd;
mem[3459] = 80'h0010d944c0550102c000;
mem[3460] = 80'h00100001ffabffabffab;
mem[3461] = 80'h0010ffcbd287edf53b94;
mem[3462] = 80'h001045a200a2557c2ff4;
mem[3463] = 80'h0010a9c2edaaa078eecc;
mem[3464] = 80'h0111c700000000000000;
mem[3465] = 80'h10100000010000010010;
mem[3466] = 80'h00109400000208004500;
mem[3467] = 80'h0010002f60350000fffd;
mem[3468] = 80'h0010d943c0550102c000;
mem[3469] = 80'h00100001ffabffabffab;
mem[3470] = 80'h0010ffcaa359c12d4256;
mem[3471] = 80'h0010fa69d225b889ffb5;
mem[3472] = 80'h0010f88ddafa00185d27;
mem[3473] = 80'h0111b600000000000000;
mem[3474] = 80'h00000000000000000000;
mem[3475] = 80'h00000000000000000000;
mem[3476] = 80'h00000000000000000000;
mem[3477] = 80'h10100000010000010010;
mem[3478] = 80'h00109400000208004500;
mem[3479] = 80'h0010002f60360000fffd;
mem[3480] = 80'h0010d942c0550102c000;
mem[3481] = 80'h00100001ffabffabffab;
mem[3482] = 80'h0010ffc9313bb445c811;
mem[3483] = 80'h00103a35a5ad8e978f06;
mem[3484] = 80'h00100a44fbde4eb56c4a;
mem[3485] = 80'h01115e00000000000000;
mem[3486] = 80'h00000000000000000000;
mem[3487] = 80'h10100000010000010010;
mem[3488] = 80'h00109400000208004500;
mem[3489] = 80'h0010002f60370000fffd;
mem[3490] = 80'h0010d941c0550102c000;
mem[3491] = 80'h00100001ffabffabffab;
mem[3492] = 80'h0010ffc840e5989db1d3;
mem[3493] = 80'h001085fe772a63625e87;
mem[3494] = 80'h00105b2aa8a3b16f2fc0;
mem[3495] = 80'h01112c00000000000000;
mem[3496] = 80'h00000000000000000000;
mem[3497] = 80'h00000000000000000000;
mem[3498] = 80'h00000000000000000000;
mem[3499] = 80'h10100000010000010010;
mem[3500] = 80'h00109400000208004500;
mem[3501] = 80'h0010002f60380000fffd;
mem[3502] = 80'h0010d940c0550102c000;
mem[3503] = 80'h00100001ffabffabffab;
mem[3504] = 80'h0010ffc778b261e7e10e;
mem[3505] = 80'h00103b447b8f56ee4c71;
mem[3506] = 80'h0010c14bab107d5c4572;
mem[3507] = 80'h0111cf00000000000000;
mem[3508] = 80'h00000000000000000000;
mem[3509] = 80'h10100000010000010010;
mem[3510] = 80'h00109400000208004500;
mem[3511] = 80'h0010002f60390000fffd;
mem[3512] = 80'h0010d93fc0550102c000;
mem[3513] = 80'h00100001ffabffabffab;
mem[3514] = 80'h0010ffc6096c4d3f98cc;
mem[3515] = 80'h0010848fa908bb1b9c77;
mem[3516] = 80'h00109090c705330c9b46;
mem[3517] = 80'h01118f00000000000000;
mem[3518] = 80'h00000000000000000000;
mem[3519] = 80'h00000000000000000000;
mem[3520] = 80'h00000000000000000000;
mem[3521] = 80'h00000000000000000000;
mem[3522] = 80'h10100000010000010010;
mem[3523] = 80'h00109400000208004500;
mem[3524] = 80'h0010002f603a0000fffd;
mem[3525] = 80'h0010d93ec0550102c000;
mem[3526] = 80'h00100001ffabffabffab;
mem[3527] = 80'h0010ffc59b0e3857128b;
mem[3528] = 80'h001044d3de808d05ecfc;
mem[3529] = 80'h001062d5da1d3f5563dd;
mem[3530] = 80'h0111ee00000000000000;
mem[3531] = 80'h10100000010000010010;
mem[3532] = 80'h00109400000208004500;
mem[3533] = 80'h0010002f603b0000fffd;
mem[3534] = 80'h0010d93dc0550102c000;
mem[3535] = 80'h00100001ffabffabffab;
mem[3536] = 80'h0010ffc4ead0148f6b49;
mem[3537] = 80'h0010fb180c0760f03c65;
mem[3538] = 80'h0010330663165ad6cc77;
mem[3539] = 80'h0111f700000000000000;
mem[3540] = 80'h00000000000000000000;
mem[3541] = 80'h00000000000000000000;
mem[3542] = 80'h00000000000000000000;
mem[3543] = 80'h10100000010000010010;
mem[3544] = 80'h00109400000208004500;
mem[3545] = 80'h0010002f603c0000fffd;
mem[3546] = 80'h0010d93cc0550102c000;
mem[3547] = 80'h00100001ffabffabffab;
mem[3548] = 80'h0010ffc3ce14fe5e7fc6;
mem[3549] = 80'h00107ba0e3160cccdd1e;
mem[3550] = 80'h0010d6979fc7f4bdadaa;
mem[3551] = 80'h0111aa00000000000000;
mem[3552] = 80'h00000000000000000000;
mem[3553] = 80'h10100000010000010010;
mem[3554] = 80'h00109400000208004500;
mem[3555] = 80'h0010002f603d0000fffd;
mem[3556] = 80'h0010d93bc0550102c000;
mem[3557] = 80'h00100001ffabffabffab;
mem[3558] = 80'h0010ffc2bfcad2860604;
mem[3559] = 80'h0010c46b3191e1390d17;
mem[3560] = 80'h0010875ccd3d2e3a7255;
mem[3561] = 80'h0111f000000000000000;
mem[3562] = 80'h00000000000000000000;
mem[3563] = 80'h00000000000000000000;
mem[3564] = 80'h00000000000000000000;
mem[3565] = 80'h10100000010000010010;
mem[3566] = 80'h00109400000208004500;
mem[3567] = 80'h0010002f603e0000fffd;
mem[3568] = 80'h0010d93ac0550102c000;
mem[3569] = 80'h00100001ffabffabffab;
mem[3570] = 80'h0010ffc12da8a7ee8c43;
mem[3571] = 80'h001004374619d7277d9c;
mem[3572] = 80'h00107519d035b9fed2d1;
mem[3573] = 80'h0111bc00000000000000;
mem[3574] = 80'h00000000000000000000;
mem[3575] = 80'h00000000000000000000;
mem[3576] = 80'h00000000000000000000;
mem[3577] = 80'h10100000010000010010;
mem[3578] = 80'h00109400000208004500;
mem[3579] = 80'h0010002f603f0000fffd;
mem[3580] = 80'h0010d939c0550102c000;
mem[3581] = 80'h00100001ffabffabffab;
mem[3582] = 80'h0010ffc05c768b36f581;
mem[3583] = 80'h0010bbfc949e3ad2ade5;
mem[3584] = 80'h001024dadbe2e8b865c5;
mem[3585] = 80'h01112900000000000000;
mem[3586] = 80'h00000000000000000000;
mem[3587] = 80'h10100000010000010010;
mem[3588] = 80'h00109400000208004500;
mem[3589] = 80'h0010002f60400000fffd;
mem[3590] = 80'h0010d938c0550102c000;
mem[3591] = 80'h00100001ffabffabffab;
mem[3592] = 80'h0010ffbfcbd386ed1e21;
mem[3593] = 80'h0010715fcc20177b09ee;
mem[3594] = 80'h001043c3a5b1467b8706;
mem[3595] = 80'h0111a700000000000000;
mem[3596] = 80'h00000000000000000000;
mem[3597] = 80'h00000000000000000000;
mem[3598] = 80'h00000000000000000000;
mem[3599] = 80'h10100000010000010010;
mem[3600] = 80'h00109400000208004500;
mem[3601] = 80'h0010002f60410000fffd;
mem[3602] = 80'h0010d937c0550102c000;
mem[3603] = 80'h00100001ffabffabffab;
mem[3604] = 80'h0010ffbeba0daa3567e3;
mem[3605] = 80'h0010ce941ea7fa8ed9a7;
mem[3606] = 80'h001012053ba3241d16c3;
mem[3607] = 80'h0111bb00000000000000;
mem[3608] = 80'h00000000000000000000;
mem[3609] = 80'h10100000010000010010;
mem[3610] = 80'h00109400000208004500;
mem[3611] = 80'h0010002f60420000fffd;
mem[3612] = 80'h0010d936c0550102c000;
mem[3613] = 80'h00100001ffabffabffab;
mem[3614] = 80'h0010ffbd286fdf5deda4;
mem[3615] = 80'h00100ec8692fcc90a96c;
mem[3616] = 80'h0010e04dea8d513c0b1a;
mem[3617] = 80'h01111f00000000000000;
mem[3618] = 80'h00000000000000000000;
mem[3619] = 80'h00000000000000000000;
mem[3620] = 80'h00000000000000000000;
mem[3621] = 80'h10100000010000010010;
mem[3622] = 80'h00109400000208004500;
mem[3623] = 80'h0010002f60430000fffd;
mem[3624] = 80'h0010d935c0550102c000;
mem[3625] = 80'h00100001ffabffabffab;
mem[3626] = 80'h0010ffbc59b1f3859466;
mem[3627] = 80'h0010b103bba821657935;
mem[3628] = 80'h0010b18807d65d8cb04a;
mem[3629] = 80'h01118700000000000000;
mem[3630] = 80'h00000000000000000000;
mem[3631] = 80'h10100000010000010010;
mem[3632] = 80'h00109400000208004500;
mem[3633] = 80'h0010002f60440000fffd;
mem[3634] = 80'h0010d934c0550102c000;
mem[3635] = 80'h00100001ffabffabffab;
mem[3636] = 80'h0010ffbb7d75195480e9;
mem[3637] = 80'h001031bb54b94d59988e;
mem[3638] = 80'h0010540faf2578f45d60;
mem[3639] = 80'h01110800000000000000;
mem[3640] = 80'h00000000000000000000;
mem[3641] = 80'h00000000000000000000;
mem[3642] = 80'h00000000000000000000;
mem[3643] = 80'h00000000000000000000;
mem[3644] = 80'h10100000010000010010;
mem[3645] = 80'h00109400000208004500;
mem[3646] = 80'h0010002f60450000fffd;
mem[3647] = 80'h0010d933c0550102c000;
mem[3648] = 80'h00100001ffabffabffab;
mem[3649] = 80'h0010ffba0cab358cf92b;
mem[3650] = 80'h00108e70863ea0ac48c7;
mem[3651] = 80'h001005c931f68eeecc86;
mem[3652] = 80'h01114100000000000000;
mem[3653] = 80'h10100000010000010010;
mem[3654] = 80'h00109400000208004500;
mem[3655] = 80'h0010002f60460000fffd;
mem[3656] = 80'h0010d932c0550102c000;
mem[3657] = 80'h00100001ffabffabffab;
mem[3658] = 80'h0010ffb99ec940e4736c;
mem[3659] = 80'h00104e2cf1b696b2380f;
mem[3660] = 80'h0010f7d4b3b1f252a401;
mem[3661] = 80'h01113c00000000000000;
mem[3662] = 80'h00000000000000000000;
mem[3663] = 80'h00000000000000000000;
mem[3664] = 80'h00000000000000000000;
mem[3665] = 80'h10100000010000010010;
mem[3666] = 80'h00109400000208004500;
mem[3667] = 80'h0010002f60470000fffd;
mem[3668] = 80'h0010d931c0550102c000;
mem[3669] = 80'h00100001ffabffabffab;
mem[3670] = 80'h0010ffb8ef176c3c0aae;
mem[3671] = 80'h0010f1e723317b47e876;
mem[3672] = 80'h0010a617b855c2ea27cb;
mem[3673] = 80'h01116700000000000000;
mem[3674] = 80'h10100000010000010010;
mem[3675] = 80'h00109400000208004500;
mem[3676] = 80'h0010002f60480000fffd;
mem[3677] = 80'h0010d930c0550102c000;
mem[3678] = 80'h00100001ffabffabffab;
mem[3679] = 80'h0010ffb7d74095465a73;
mem[3680] = 80'h00104f5d2f944ecbfa88;
mem[3681] = 80'h00103cff1209219082e5;
mem[3682] = 80'h01115c00000000000000;
mem[3683] = 80'h00000000000000000000;
mem[3684] = 80'h00000000000000000000;
mem[3685] = 80'h00000000000000000000;
mem[3686] = 80'h10100000010000010010;
mem[3687] = 80'h00109400000208004500;
mem[3688] = 80'h0010002f60490000fffd;
mem[3689] = 80'h0010d92fc0550102c000;
mem[3690] = 80'h00100001ffabffabffab;
mem[3691] = 80'h0010ffb6a69eb99e23b1;
mem[3692] = 80'h0010f096fd13a33e2b01;
mem[3693] = 80'h00106d18e8576a6857d0;
mem[3694] = 80'h01115f00000000000000;
mem[3695] = 80'h00000000000000000000;
mem[3696] = 80'h10100000010000010010;
mem[3697] = 80'h00109400000208004500;
mem[3698] = 80'h0010002f604a0000fffd;
mem[3699] = 80'h0010d92ec0550102c000;
mem[3700] = 80'h00100001ffabffabffab;
mem[3701] = 80'h0010ffb534fcccf6a9f6;
mem[3702] = 80'h001030ca8a9b95205b8a;
mem[3703] = 80'h00109f5df5f212e1ca48;
mem[3704] = 80'h01113800000000000000;
mem[3705] = 80'h00000000000000000000;
mem[3706] = 80'h00000000000000000000;
mem[3707] = 80'h00000000000000000000;
mem[3708] = 80'h00000000000000000000;
mem[3709] = 80'h10100000010000010010;
mem[3710] = 80'h00109400000208004500;
mem[3711] = 80'h0010002f604b0000fffd;
mem[3712] = 80'h0010d92dc0550102c000;
mem[3713] = 80'h00100001ffabffabffab;
mem[3714] = 80'h0010ffb44522e02ed034;
mem[3715] = 80'h00108f01581c78d58b93;
mem[3716] = 80'h0010ce95d4a87b52685c;
mem[3717] = 80'h0111e100000000000000;
mem[3718] = 80'h00000000000000000000;
mem[3719] = 80'h10100000010000010010;
mem[3720] = 80'h00109400000208004500;
mem[3721] = 80'h0010002f604c0000fffd;
mem[3722] = 80'h0010d92cc0550102c000;
mem[3723] = 80'h00100001ffabffabffab;
mem[3724] = 80'h0010ffb361e60affc4bb;
mem[3725] = 80'h00100fb9b70d14e96ae9;
mem[3726] = 80'h00102b3719db42f8dab0;
mem[3727] = 80'h01114200000000000000;
mem[3728] = 80'h00000000000000000000;
mem[3729] = 80'h00000000000000000000;
mem[3730] = 80'h00000000000000000000;
mem[3731] = 80'h10100000010000010010;
mem[3732] = 80'h00109400000208004500;
mem[3733] = 80'h0010002f604d0000fffd;
mem[3734] = 80'h0010d92bc0550102c000;
mem[3735] = 80'h00100001ffabffabffab;
mem[3736] = 80'h0010ffb210382627bd79;
mem[3737] = 80'h0010b072658af91cba60;
mem[3738] = 80'h00107ae7d311f4f133a5;
mem[3739] = 80'h0111e900000000000000;
mem[3740] = 80'h00000000000000000000;
mem[3741] = 80'h10100000010000010010;
mem[3742] = 80'h00109400000208004500;
mem[3743] = 80'h0010002f604e0000fffd;
mem[3744] = 80'h0010d92ac0550102c000;
mem[3745] = 80'h00100001ffabffabffab;
mem[3746] = 80'h0010ffb1825a534f373e;
mem[3747] = 80'h0010702e1202cf02caeb;
mem[3748] = 80'h001088a2cea47f8f1f4b;
mem[3749] = 80'h0111e000000000000000;
mem[3750] = 80'h00000000000000000000;
mem[3751] = 80'h10100000010000010010;
mem[3752] = 80'h00109400000208004500;
mem[3753] = 80'h0010002f604f0000fffd;
mem[3754] = 80'h0010d929c0550102c000;
mem[3755] = 80'h00100001ffabffabffab;
mem[3756] = 80'h0010ffb0f3847f974efc;
mem[3757] = 80'h0010cfe5c08522f71a92;
mem[3758] = 80'h0010d961c5dfd03784e8;
mem[3759] = 80'h01112d00000000000000;
mem[3760] = 80'h00000000000000000000;
mem[3761] = 80'h00000000000000000000;
mem[3762] = 80'h00000000000000000000;
mem[3763] = 80'h10100000010000010010;
mem[3764] = 80'h00109400000208004500;
mem[3765] = 80'h0010002f60500000fffd;
mem[3766] = 80'h0010d928c0550102c000;
mem[3767] = 80'h00100001ffabffabffab;
mem[3768] = 80'h0010ffaff2f5a1bb9685;
mem[3769] = 80'h00100d5a0b48a41aef26;
mem[3770] = 80'h0010bc662ecf3db182b2;
mem[3771] = 80'h01116700000000000000;
mem[3772] = 80'h00000000000000000000;
mem[3773] = 80'h10100000010000010010;
mem[3774] = 80'h00109400000208004500;
mem[3775] = 80'h0010002f60510000fffd;
mem[3776] = 80'h0010d927c0550102c000;
mem[3777] = 80'h00100001ffabffabffab;
mem[3778] = 80'h0010ffae832b8d63ef47;
mem[3779] = 80'h0010b291d9cf49ef3f6f;
mem[3780] = 80'h0010eda0b0194c43405f;
mem[3781] = 80'h01115000000000000000;
mem[3782] = 80'h00000000000000000000;
mem[3783] = 80'h00000000000000000000;
mem[3784] = 80'h00000000000000000000;
mem[3785] = 80'h10100000010000010010;
mem[3786] = 80'h00109400000208004500;
mem[3787] = 80'h0010002f60520000fffd;
mem[3788] = 80'h0010d926c0550102c000;
mem[3789] = 80'h00100001ffabffabffab;
mem[3790] = 80'h0010ffad1149f80b6500;
mem[3791] = 80'h001072cdae477ff14823;
mem[3792] = 80'h00101feffee3896f3339;
mem[3793] = 80'h01117700000000000000;
mem[3794] = 80'h00000000000000000000;
mem[3795] = 80'h10100000010000010010;
mem[3796] = 80'h00109400000208004500;
mem[3797] = 80'h0010002f60530000fffd;
mem[3798] = 80'h0010d925c0550102c000;
mem[3799] = 80'h00100001ffabffabffab;
mem[3800] = 80'h0010ffac6097d4d31cc2;
mem[3801] = 80'h0010cd067cc092049862;
mem[3802] = 80'h00104ea0c9572142664b;
mem[3803] = 80'h01110a00000000000000;
mem[3804] = 80'h00000000000000000000;
mem[3805] = 80'h00000000000000000000;
mem[3806] = 80'h00000000000000000000;
mem[3807] = 80'h00000000000000000000;
mem[3808] = 80'h10100000010000010010;
mem[3809] = 80'h00109400000208004500;
mem[3810] = 80'h0010002f60540000fffd;
mem[3811] = 80'h0010d924c0550102c000;
mem[3812] = 80'h00100001ffabffabffab;
mem[3813] = 80'h0010ffab44533e02084d;
mem[3814] = 80'h00104dbe93d1fe387941;
mem[3815] = 80'h0010abb623f14cc8a07d;
mem[3816] = 80'h0111bd00000000000000;
mem[3817] = 80'h10100000010000010010;
mem[3818] = 80'h00109400000208004500;
mem[3819] = 80'h0010002f60550000fffd;
mem[3820] = 80'h0010d923c0550102c000;
mem[3821] = 80'h00100001ffabffabffab;
mem[3822] = 80'h0010ffaa358d12da718f;
mem[3823] = 80'h0010f275415613cda900;
mem[3824] = 80'h0010faf914cb45c98b8e;
mem[3825] = 80'h0111fc00000000000000;
mem[3826] = 80'h00000000000000000000;
mem[3827] = 80'h00000000000000000000;
mem[3828] = 80'h00000000000000000000;
mem[3829] = 80'h10100000010000010010;
mem[3830] = 80'h00109400000208004500;
mem[3831] = 80'h0010002f60560000fffd;
mem[3832] = 80'h0010d922c0550102c000;
mem[3833] = 80'h00100001ffabffabffab;
mem[3834] = 80'h0010ffa9a7ef67b2fbc8;
mem[3835] = 80'h0010322936de25d3d943;
mem[3836] = 80'h00100823f4a98fc10846;
mem[3837] = 80'h01119f00000000000000;
mem[3838] = 80'h00000000000000000000;
mem[3839] = 80'h10100000010000010010;
mem[3840] = 80'h00109400000208004500;
mem[3841] = 80'h0010002f60570000fffd;
mem[3842] = 80'h0010d921c0550102c000;
mem[3843] = 80'h00100001ffabffabffab;
mem[3844] = 80'h0010ffa8d6314b6a820a;
mem[3845] = 80'h00108de2e459c8260902;
mem[3846] = 80'h0010596cc3defb9e4786;
mem[3847] = 80'h01118d00000000000000;
mem[3848] = 80'h00000000000000000000;
mem[3849] = 80'h00000000000000000000;
mem[3850] = 80'h00000000000000000000;
mem[3851] = 80'h10100000010000010010;
mem[3852] = 80'h00109400000208004500;
mem[3853] = 80'h0010002f60580000fffd;
mem[3854] = 80'h0010d920c0550102c000;
mem[3855] = 80'h00100001ffabffabffab;
mem[3856] = 80'h0010ffa7ee66b210d2d7;
mem[3857] = 80'h00103358e8fcfdaa1bc4;
mem[3858] = 80'h0010c308553c3e987434;
mem[3859] = 80'h01117c00000000000000;
mem[3860] = 80'h00000000000000000000;
mem[3861] = 80'h10100000010000010010;
mem[3862] = 80'h00109400000208004500;
mem[3863] = 80'h0010002f60590000fffd;
mem[3864] = 80'h0010d91fc0550102c000;
mem[3865] = 80'h00100001ffabffabffab;
mem[3866] = 80'h0010ffa69fb89ec8ab15;
mem[3867] = 80'h00108c933a7b105fcbc4;
mem[3868] = 80'h001092799f1641923e9d;
mem[3869] = 80'h01112f00000000000000;
mem[3870] = 80'h00000000000000000000;
mem[3871] = 80'h00000000000000000000;
mem[3872] = 80'h00000000000000000000;
mem[3873] = 80'h00000000000000000000;
mem[3874] = 80'h10100000010000010010;
mem[3875] = 80'h00109400000208004500;
mem[3876] = 80'h0010002f605a0000fffd;
mem[3877] = 80'h0010d91ec0550102c000;
mem[3878] = 80'h00100001ffabffabffab;
mem[3879] = 80'h0010ffa50ddaeba02152;
mem[3880] = 80'h00104ccf4df32641bb47;
mem[3881] = 80'h001060b52b8cdce38210;
mem[3882] = 80'h01116a00000000000000;
mem[3883] = 80'h10100000010000010010;
mem[3884] = 80'h00109400000208004500;
mem[3885] = 80'h0010002f605b0000fffd;
mem[3886] = 80'h0010d91dc0550102c000;
mem[3887] = 80'h00100001ffabffabffab;
mem[3888] = 80'h0010ffa47c04c7785890;
mem[3889] = 80'h0010f3049f74cbb46ac6;
mem[3890] = 80'h001031db787df0109576;
mem[3891] = 80'h01119000000000000000;
mem[3892] = 80'h00000000000000000000;
mem[3893] = 80'h00000000000000000000;
mem[3894] = 80'h00000000000000000000;
mem[3895] = 80'h10100000010000010010;
mem[3896] = 80'h00109400000208004500;
mem[3897] = 80'h0010002f605c0000fffd;
mem[3898] = 80'h0010d91cc0550102c000;
mem[3899] = 80'h00100001ffabffabffab;
mem[3900] = 80'h0010ffa358c02da94c1f;
mem[3901] = 80'h001073bc7065a7888ba5;
mem[3902] = 80'h0010d4c05ec2e2ba2b7d;
mem[3903] = 80'h01111900000000000000;
mem[3904] = 80'h00000000000000000000;
mem[3905] = 80'h10100000010000010010;
mem[3906] = 80'h00109400000208004500;
mem[3907] = 80'h0010002f605d0000fffd;
mem[3908] = 80'h0010d91bc0550102c000;
mem[3909] = 80'h00100001ffabffabffab;
mem[3910] = 80'h0010ffa2291e017135dd;
mem[3911] = 80'h0010cc77a2e24a7d5ba4;
mem[3912] = 80'h00108582a5f25ea712ed;
mem[3913] = 80'h01117c00000000000000;
mem[3914] = 80'h00000000000000000000;
mem[3915] = 80'h00000000000000000000;
mem[3916] = 80'h00000000000000000000;
mem[3917] = 80'h10100000010000010010;
mem[3918] = 80'h00109400000208004500;
mem[3919] = 80'h0010002f605e0000fffd;
mem[3920] = 80'h0010d91ac0550102c000;
mem[3921] = 80'h00100001ffabffabffab;
mem[3922] = 80'h0010ffa1bb7c7419bf9a;
mem[3923] = 80'h00100c2bd56a7c632b27;
mem[3924] = 80'h0010774e11befe5e806a;
mem[3925] = 80'h0111b600000000000000;
mem[3926] = 80'h00000000000000000000;
mem[3927] = 80'h00000000000000000000;
mem[3928] = 80'h00000000000000000000;
mem[3929] = 80'h10100000010000010010;
mem[3930] = 80'h00109400000208004500;
mem[3931] = 80'h0010002f605f0000fffd;
mem[3932] = 80'h0010d919c0550102c000;
mem[3933] = 80'h00100001ffabffabffab;
mem[3934] = 80'h0010ffa0caa258c1c658;
mem[3935] = 80'h0010b3e007ed9196fba5;
mem[3936] = 80'h0010264221568509c95e;
mem[3937] = 80'h0111d900000000000000;
mem[3938] = 80'h00000000000000000000;
mem[3939] = 80'h10100000010000010010;
mem[3940] = 80'h00109400000208004500;
mem[3941] = 80'h0010002f60600000fffd;
mem[3942] = 80'h0010d918c0550102c000;
mem[3943] = 80'h00100001ffabffabffab;
mem[3944] = 80'h0010ff9fb99fc8400f69;
mem[3945] = 80'h0010895442f171b8c07c;
mem[3946] = 80'h0010bd11018ab1cb6e8b;
mem[3947] = 80'h01113500000000000000;
mem[3948] = 80'h00000000000000000000;
mem[3949] = 80'h00000000000000000000;
mem[3950] = 80'h00000000000000000000;
mem[3951] = 80'h10100000010000010010;
mem[3952] = 80'h00109400000208004500;
mem[3953] = 80'h0010002f60610000fffd;
mem[3954] = 80'h0010d917c0550102c000;
mem[3955] = 80'h00100001ffabffabffab;
mem[3956] = 80'h0010ff9ec841e49876ab;
mem[3957] = 80'h0010369f90769c4d103d;
mem[3958] = 80'h0010ec5e36dc45ee5e9c;
mem[3959] = 80'h01110e00000000000000;
mem[3960] = 80'h00000000000000000000;
mem[3961] = 80'h10100000010000010010;
mem[3962] = 80'h00109400000208004500;
mem[3963] = 80'h0010002f60620000fffd;
mem[3964] = 80'h0010d916c0550102c000;
mem[3965] = 80'h00100001ffabffabffab;
mem[3966] = 80'h0010ff9d5a2391f0fcec;
mem[3967] = 80'h0010f6c3e7feaa5360fe;
mem[3968] = 80'h00101e9f4eadbfd681ca;
mem[3969] = 80'h01114000000000000000;
mem[3970] = 80'h00000000000000000000;
mem[3971] = 80'h00000000000000000000;
mem[3972] = 80'h00000000000000000000;
mem[3973] = 80'h10100000010000010010;
mem[3974] = 80'h00109400000208004500;
mem[3975] = 80'h0010002f60630000fffd;
mem[3976] = 80'h0010d915c0550102c000;
mem[3977] = 80'h00100001ffabffabffab;
mem[3978] = 80'h0010ff9c2bfdbd28852e;
mem[3979] = 80'h00104908357947a6b0bf;
mem[3980] = 80'h00104fd0795751d552fd;
mem[3981] = 80'h0111cc00000000000000;
mem[3982] = 80'h00000000000000000000;
mem[3983] = 80'h10100000010000010010;
mem[3984] = 80'h00109400000208004500;
mem[3985] = 80'h0010002f60640000fffd;
mem[3986] = 80'h0010d914c0550102c000;
mem[3987] = 80'h00100001ffabffabffab;
mem[3988] = 80'h0010ff9b0f3957f991a1;
mem[3989] = 80'h0010c9b0da682b9a521c;
mem[3990] = 80'h0010aa845b3bdf524124;
mem[3991] = 80'h0111f200000000000000;
mem[3992] = 80'h00000000000000000000;
mem[3993] = 80'h00000000000000000000;
mem[3994] = 80'h00000000000000000000;
mem[3995] = 80'h00000000000000000000;
mem[3996] = 80'h10100000010000010010;
mem[3997] = 80'h00109400000208004500;
mem[3998] = 80'h0010002f60650000fffd;
mem[3999] = 80'h0010d913c0550102c000;
mem[4000] = 80'h00100001ffabffabffab;
mem[4001] = 80'h0010ff9a7ee77b21e863;
mem[4002] = 80'h0010767b08efc66f825c;
mem[4003] = 80'h0010fbf85dc8fb6c515b;
mem[4004] = 80'h0111e000000000000000;
mem[4005] = 80'h10100000010000010010;
mem[4006] = 80'h00109400000208004500;
mem[4007] = 80'h0010002f60660000fffd;
mem[4008] = 80'h0010d912c0550102c000;
mem[4009] = 80'h00100001ffabffabffab;
mem[4010] = 80'h0010ff99ec850e496224;
mem[4011] = 80'h0010b6277f67f071f29f;
mem[4012] = 80'h0010093925995b1c1237;
mem[4013] = 80'h0111b000000000000000;
mem[4014] = 80'h00000000000000000000;
mem[4015] = 80'h00000000000000000000;
mem[4016] = 80'h00000000000000000000;
mem[4017] = 80'h10100000010000010010;
mem[4018] = 80'h00109400000208004500;
mem[4019] = 80'h0010002f60670000fffd;
mem[4020] = 80'h0010d911c0550102c000;
mem[4021] = 80'h00100001ffabffabffab;
mem[4022] = 80'h0010ff989d5b22911be6;
mem[4023] = 80'h001009ecade01d8422de;
mem[4024] = 80'h0010587612efc0eb9359;
mem[4025] = 80'h01118b00000000000000;
mem[4026] = 80'h10100000010000010010;
mem[4027] = 80'h00109400000208004500;
mem[4028] = 80'h0010002f60680000fffd;
mem[4029] = 80'h0010d910c0550102c000;
mem[4030] = 80'h00100001ffabffabffab;
mem[4031] = 80'h0010ff97a50cdbeb4b3b;
mem[4032] = 80'h0010b756a14528083018;
mem[4033] = 80'h0010c21284653c4ac9ca;
mem[4034] = 80'h01118800000000000000;
mem[4035] = 80'h00000000000000000000;
mem[4036] = 80'h00000000000000000000;
mem[4037] = 80'h00000000000000000000;
mem[4038] = 80'h10100000010000010010;
mem[4039] = 80'h00109400000208004500;
mem[4040] = 80'h0010002f60690000fffd;
mem[4041] = 80'h0010d90fc0550102c000;
mem[4042] = 80'h00100001ffabffabffab;
mem[4043] = 80'h0010ff96d4d2f73332f9;
mem[4044] = 80'h0010089d73c2c5fde099;
mem[4045] = 80'h0010934be72663dc9702;
mem[4046] = 80'h01112b00000000000000;
mem[4047] = 80'h00000000000000000000;
mem[4048] = 80'h10100000010000010010;
mem[4049] = 80'h00109400000208004500;
mem[4050] = 80'h0010002f606a0000fffd;
mem[4051] = 80'h0010d90ec0550102c000;
mem[4052] = 80'h00100001ffabffabffab;
mem[4053] = 80'h0010ff9546b0825bb8be;
mem[4054] = 80'h0010c8c1044af3e3901a;
mem[4055] = 80'h00106187530e7882c1a7;
mem[4056] = 80'h0111bc00000000000000;
mem[4057] = 80'h00000000000000000000;
mem[4058] = 80'h00000000000000000000;
mem[4059] = 80'h00000000000000000000;
mem[4060] = 80'h10100000010000010010;
mem[4061] = 80'h00109400000208004500;
mem[4062] = 80'h0010002f606b0000fffd;
mem[4063] = 80'h0010d90dc0550102c000;
mem[4064] = 80'h00100001ffabffabffab;
mem[4065] = 80'h0010ff94376eae83c17c;
mem[4066] = 80'h0010770ad6cd1e16401c;
mem[4067] = 80'h0010305c3f963c24dcce;
mem[4068] = 80'h01111100000000000000;
mem[4069] = 80'h00000000000000000000;
mem[4070] = 80'h10100000010000010010;
mem[4071] = 80'h00109400000208004500;
mem[4072] = 80'h0010002f606c0000fffd;
mem[4073] = 80'h0010d90cc0550102c000;
mem[4074] = 80'h00100001ffabffabffab;
mem[4075] = 80'h0010ff9313aa4452d5f3;
mem[4076] = 80'h0010f7b239dc722aa167;
mem[4077] = 80'h0010d5cdc38cf304e2a8;
mem[4078] = 80'h01115e00000000000000;
mem[4079] = 80'h00000000000000000000;
mem[4080] = 80'h00000000000000000000;
mem[4081] = 80'h00000000000000000000;
mem[4082] = 80'h10100000010000010010;
mem[4083] = 80'h00109400000208004500;
mem[4084] = 80'h0010002f606d0000fffd;
mem[4085] = 80'h0010d90bc0550102c000;
mem[4086] = 80'h00100001ffabffabffab;
mem[4087] = 80'h0010ff926274688aac31;
mem[4088] = 80'h00104879eb5b9fdf70fe;
mem[4089] = 80'h001084294a6075c5ed8e;
mem[4090] = 80'h0111b800000000000000;
mem[4091] = 80'h00000000000000000000;
mem[4092] = 80'h10100000010000010010;
mem[4093] = 80'h00109400000208004500;
mem[4094] = 80'h0010002f606e0000fffd;
mem[4095] = 80'h0010d90ac0550102c000;
mem[4096] = 80'h00100001ffabffabffab;
mem[4097] = 80'h0010ff91f0161de22676;
mem[4098] = 80'h001088259cd3a9c10075;
mem[4099] = 80'h0010766c57632e511a2c;
mem[4100] = 80'h01118500000000000000;
mem[4101] = 80'h00000000000000000000;
mem[4102] = 80'h00000000000000000000;
mem[4103] = 80'h00000000000000000000;
mem[4104] = 80'h10100000010000010010;
mem[4105] = 80'h00109400000208004500;
mem[4106] = 80'h0010002f606f0000fffd;
mem[4107] = 80'h0010d909c0550102c000;
mem[4108] = 80'h00100001ffabffabffab;
mem[4109] = 80'h0010ff9081c8313a5fb4;
mem[4110] = 80'h001037ee4e544434d07c;
mem[4111] = 80'h001027a7051e258f7195;
mem[4112] = 80'h01116200000000000000;
mem[4113] = 80'h00000000000000000000;
mem[4114] = 80'h10100000010000010010;
mem[4115] = 80'h00109400000208004500;
mem[4116] = 80'h0010002f60700000fffd;
mem[4117] = 80'h0010d908c0550102c000;
mem[4118] = 80'h00100001ffabffabffab;
mem[4119] = 80'h0010ff8f80b9ef1687cd;
mem[4120] = 80'h0010f5518599c2d92588;
mem[4121] = 80'h001042ad22d83fbacff3;
mem[4122] = 80'h0111b900000000000000;
mem[4123] = 80'h00000000000000000000;
mem[4124] = 80'h00000000000000000000;
mem[4125] = 80'h00000000000000000000;
mem[4126] = 80'h10100000010000010010;
mem[4127] = 80'h00109400000208004500;
mem[4128] = 80'h0010002f60710000fffd;
mem[4129] = 80'h0010d907c0550102c000;
mem[4130] = 80'h00100001ffabffabffab;
mem[4131] = 80'h0010ff8ef167c3cefe0f;
mem[4132] = 80'h00104a9a571e2f2cf5f1;
mem[4133] = 80'h0010136e29e6481d5ca6;
mem[4134] = 80'h01113900000000000000;
mem[4135] = 80'h00000000000000000000;
mem[4136] = 80'h10100000010000010010;
mem[4137] = 80'h00109400000208004500;
mem[4138] = 80'h0010002f60720000fffd;
mem[4139] = 80'h0010d906c0550102c000;
mem[4140] = 80'h00100001ffabffabffab;
mem[4141] = 80'h0010ff8d6305b6a67448;
mem[4142] = 80'h00108ac62096193285bb;
mem[4143] = 80'h0010e10e5124f51d91c8;
mem[4144] = 80'h01119c00000000000000;
mem[4145] = 80'h00000000000000000000;
mem[4146] = 80'h00000000000000000000;
mem[4147] = 80'h00000000000000000000;
mem[4148] = 80'h10100000010000010010;
mem[4149] = 80'h00109400000208004500;
mem[4150] = 80'h0010002f60730000fffd;
mem[4151] = 80'h0010d905c0550102c000;
mem[4152] = 80'h00100001ffabffabffab;
mem[4153] = 80'h0010ff8c12db9a7e0d8a;
mem[4154] = 80'h0010350df211f4c755f2;
mem[4155] = 80'h0010b0c8cfed5229c33f;
mem[4156] = 80'h01114100000000000000;
mem[4157] = 80'h00000000000000000000;
mem[4158] = 80'h10100000010000010010;
mem[4159] = 80'h00109400000208004500;
mem[4160] = 80'h0010002f60740000fffd;
mem[4161] = 80'h0010d904c0550102c000;
mem[4162] = 80'h00100001ffabffabffab;
mem[4163] = 80'h0010ff8b361f70af1905;
mem[4164] = 80'h0010b5b51d0098fbb4c9;
mem[4165] = 80'h00105554ffd0caae3614;
mem[4166] = 80'h01114400000000000000;
mem[4167] = 80'h00000000000000000000;
mem[4168] = 80'h00000000000000000000;
mem[4169] = 80'h00000000000000000000;
mem[4170] = 80'h10100000010000010010;
mem[4171] = 80'h00109400000208004500;
mem[4172] = 80'h0010002f60750000fffd;
mem[4173] = 80'h0010d903c0550102c000;
mem[4174] = 80'h00100001ffabffabffab;
mem[4175] = 80'h0010ff8a47c15c7760c7;
mem[4176] = 80'h00100a7ecf87750e6490;
mem[4177] = 80'h00100491124030258cc4;
mem[4178] = 80'h01119800000000000000;
mem[4179] = 80'h00000000000000000000;
mem[4180] = 80'h10100000010000010010;
mem[4181] = 80'h00109400000208004500;
mem[4182] = 80'h0010002f60760000fffd;
mem[4183] = 80'h0010d902c0550102c000;
mem[4184] = 80'h00100001ffabffabffab;
mem[4185] = 80'h0010ff89d5a3291fea80;
mem[4186] = 80'h0010ca22b80f43102bdb;
mem[4187] = 80'h0010f62bcfe85f98b148;
mem[4188] = 80'h0111c900000000000000;
mem[4189] = 80'h00000000000000000000;
mem[4190] = 80'h00000000000000000000;
mem[4191] = 80'h00000000000000000000;
mem[4192] = 80'h10100000010000010010;
mem[4193] = 80'h00109400000208004500;
mem[4194] = 80'h0010002f60770000fffd;
mem[4195] = 80'h0010d901c0550102c000;
mem[4196] = 80'h00100001ffabffabffab;
mem[4197] = 80'h0010ff88a47d05c79342;
mem[4198] = 80'h001075e96a88aee5fb92;
mem[4199] = 80'h0010a7ed51183e93093c;
mem[4200] = 80'h01116800000000000000;
mem[4201] = 80'h00000000000000000000;
mem[4202] = 80'h10100000010000010010;
mem[4203] = 80'h00109400000208004500;
mem[4204] = 80'h0010002f60780000fffd;
mem[4205] = 80'h0010d900c0550102c000;
mem[4206] = 80'h00100001ffabffabffab;
mem[4207] = 80'h0010ff879c2afcbdc39f;
mem[4208] = 80'h0010cb53662d9b69e92f;
mem[4209] = 80'h00103d5d64784b2543b7;
mem[4210] = 80'h01114800000000000000;
mem[4211] = 80'h00000000000000000000;
mem[4212] = 80'h00000000000000000000;
mem[4213] = 80'h00000000000000000000;
mem[4214] = 80'h00000000000000000000;
mem[4215] = 80'h10100000010000010010;
mem[4216] = 80'h00109400000208004500;
mem[4217] = 80'h0010002f60790000fffd;
mem[4218] = 80'h0010d8ffc0550102c000;
mem[4219] = 80'h00100001ffabffabffab;
mem[4220] = 80'h0010ff86edf4d065ba5d;
mem[4221] = 80'h00107498b4aa769c3956;
mem[4222] = 80'h00106c9e6fecd18823db;
mem[4223] = 80'h01116e00000000000000;
mem[4224] = 80'h00000000000000000000;
mem[4225] = 80'h10100000010000010010;
mem[4226] = 80'h00109400000208004500;
mem[4227] = 80'h0010002f607a0000fffd;
mem[4228] = 80'h0010d8fec0550102c000;
mem[4229] = 80'h00100001ffabffabffab;
mem[4230] = 80'h0010ff857f96a50d301a;
mem[4231] = 80'h0010b4c4c322408249dd;
mem[4232] = 80'h00109edb729997b5661a;
mem[4233] = 80'h01114900000000000000;
mem[4234] = 80'h00000000000000000000;
mem[4235] = 80'h00000000000000000000;
mem[4236] = 80'h00000000000000000000;
mem[4237] = 80'h10100000010000010010;
mem[4238] = 80'h00109400000208004500;
mem[4239] = 80'h0010002f607b0000fffd;
mem[4240] = 80'h0010d8fdc0550102c000;
mem[4241] = 80'h00100001ffabffabffab;
mem[4242] = 80'h0010ff840e4889d549d8;
mem[4243] = 80'h00100b0f11a5ad779954;
mem[4244] = 80'h0010cf0bb8f93296c209;
mem[4245] = 80'h01110a00000000000000;
mem[4246] = 80'h00000000000000000000;
mem[4247] = 80'h10100000010000010010;
mem[4248] = 80'h00109400000208004500;
mem[4249] = 80'h0010002f607c0000fffd;
mem[4250] = 80'h0010d8fcc0550102c000;
mem[4251] = 80'h00100001ffabffabffab;
mem[4252] = 80'h0010ff832a8c63045d57;
mem[4253] = 80'h00108bb7feb4c14b782f;
mem[4254] = 80'h00102a9a4412e2bf21c0;
mem[4255] = 80'h0111c500000000000000;
mem[4256] = 80'h00000000000000000000;
mem[4257] = 80'h00000000000000000000;
mem[4258] = 80'h00000000000000000000;
mem[4259] = 80'h10100000010000010010;
mem[4260] = 80'h00109400000208004500;
mem[4261] = 80'h0010002f607d0000fffd;
mem[4262] = 80'h0010d8fbc0550102c000;
mem[4263] = 80'h00100001ffabffabffab;
mem[4264] = 80'h0010ff825b524fdc2495;
mem[4265] = 80'h0010347c2c332cbea836;
mem[4266] = 80'h00107b5265c3197368f2;
mem[4267] = 80'h0111e200000000000000;
mem[4268] = 80'h00000000000000000000;
mem[4269] = 80'h10100000010000010010;
mem[4270] = 80'h00109400000208004500;
mem[4271] = 80'h0010002f607e0000fffd;
mem[4272] = 80'h0010d8fac0550102c000;
mem[4273] = 80'h00100001ffabffabffab;
mem[4274] = 80'h0010ff81c9303ab4aed2;
mem[4275] = 80'h0010f4205bbb1aa0d8bc;
mem[4276] = 80'h00108924496937b91691;
mem[4277] = 80'h01118c00000000000000;
mem[4278] = 80'h00000000000000000000;
mem[4279] = 80'h00000000000000000000;
mem[4280] = 80'h00000000000000000000;
mem[4281] = 80'h10100000010000010010;
mem[4282] = 80'h00109400000208004500;
mem[4283] = 80'h0010002f607f0000fffd;
mem[4284] = 80'h0010d8f9c0550102c000;
mem[4285] = 80'h00100001ffabffabffab;
mem[4286] = 80'h0010ff80b8ee166cd710;
mem[4287] = 80'h00104beb893cf7550935;
mem[4288] = 80'h0010d8c3b39cf72e778c;
mem[4289] = 80'h01111100000000000000;
mem[4290] = 80'h00000000000000000000;
mem[4291] = 80'h10100000010000010010;
mem[4292] = 80'h00109400000208004500;
mem[4293] = 80'h0010002f60800000fffd;
mem[4294] = 80'h0010d8f8c0550102c000;
mem[4295] = 80'h00100001ffabffabffab;
mem[4296] = 80'h0010ff7f97a40ddb0051;
mem[4297] = 80'h0010dead3841ac0646cd;
mem[4298] = 80'h00101712e3da55a123a0;
mem[4299] = 80'h0111f000000000000000;
mem[4300] = 80'h00000000000000000000;
mem[4301] = 80'h00000000000000000000;
mem[4302] = 80'h00000000000000000000;
mem[4303] = 80'h10100000010000010010;
mem[4304] = 80'h00109400000208004500;
mem[4305] = 80'h0010002f60810000fffd;
mem[4306] = 80'h0010d8f7c0550102c000;
mem[4307] = 80'h00100001ffabffabffab;
mem[4308] = 80'h0010ff7ee67a21037993;
mem[4309] = 80'h00106166eac641f396b4;
mem[4310] = 80'h001046d1e8c92adb6204;
mem[4311] = 80'h01115e00000000000000;
mem[4312] = 80'h00000000000000000000;
mem[4313] = 80'h10100000010000010010;
mem[4314] = 80'h00109400000208004500;
mem[4315] = 80'h0010002f60820000fffd;
mem[4316] = 80'h0010d8f6c0550102c000;
mem[4317] = 80'h00100001ffabffabffab;
mem[4318] = 80'h0010ff7d7418546bf3d4;
mem[4319] = 80'h0010a13a9d4e77ede67f;
mem[4320] = 80'h0010b4993999b8595c0f;
mem[4321] = 80'h01117500000000000000;
mem[4322] = 80'h00000000000000000000;
mem[4323] = 80'h00000000000000000000;
mem[4324] = 80'h00000000000000000000;
mem[4325] = 80'h10100000010000010010;
mem[4326] = 80'h00109400000208004500;
mem[4327] = 80'h0010002f60830000fffd;
mem[4328] = 80'h0010d8f5c0550102c000;
mem[4329] = 80'h00100001ffabffabffab;
mem[4330] = 80'h0010ff7c05c678b38a16;
mem[4331] = 80'h00101ef14fc99a183636;
mem[4332] = 80'h0010e55fa78a2b4dd79b;
mem[4333] = 80'h0111f200000000000000;
mem[4334] = 80'h00000000000000000000;
mem[4335] = 80'h10100000010000010010;
mem[4336] = 80'h00109400000208004500;
mem[4337] = 80'h0010002f60840000fffd;
mem[4338] = 80'h0010d8f4c0550102c000;
mem[4339] = 80'h00100001ffabffabffab;
mem[4340] = 80'h0010ff7b210292629e99;
mem[4341] = 80'h00109e49a0d8f624d78a;
mem[4342] = 80'h0010004198730869472c;
mem[4343] = 80'h01114b00000000000000;
mem[4344] = 80'h00000000000000000000;
mem[4345] = 80'h00000000000000000000;
mem[4346] = 80'h00000000000000000000;
mem[4347] = 80'h10100000010000010010;
mem[4348] = 80'h00109400000208004500;
mem[4349] = 80'h0010002f60850000fffd;
mem[4350] = 80'h0010d8f3c0550102c000;
mem[4351] = 80'h00100001ffabffabffab;
mem[4352] = 80'h0010ff7a50dcbebae75b;
mem[4353] = 80'h00102182725f1bd107cb;
mem[4354] = 80'h0010510eaf0651566e55;
mem[4355] = 80'h01111600000000000000;
mem[4356] = 80'h00000000000000000000;
mem[4357] = 80'h10100000010000010010;
mem[4358] = 80'h00109400000208004500;
mem[4359] = 80'h0010002f60860000fffd;
mem[4360] = 80'h0010d8f2c0550102c000;
mem[4361] = 80'h00100001ffabffabffab;
mem[4362] = 80'h0010ff79c2becbd26d1c;
mem[4363] = 80'h0010e1de05d72dcf7718;
mem[4364] = 80'h0010a3cca46e2f332402;
mem[4365] = 80'h01116e00000000000000;
mem[4366] = 80'h00000000000000000000;
mem[4367] = 80'h00000000000000000000;
mem[4368] = 80'h00000000000000000000;
mem[4369] = 80'h10100000010000010010;
mem[4370] = 80'h00109400000208004500;
mem[4371] = 80'h0010002f60870000fffd;
mem[4372] = 80'h0010d8f1c0550102c000;
mem[4373] = 80'h00100001ffabffabffab;
mem[4374] = 80'h0010ff78b360e70a14de;
mem[4375] = 80'h00105e15d750c03aa759;
mem[4376] = 80'h0010f28393bf2d0aa4f9;
mem[4377] = 80'h01113d00000000000000;
mem[4378] = 80'h00000000000000000000;
mem[4379] = 80'h10100000010000010010;
mem[4380] = 80'h00109400000208004500;
mem[4381] = 80'h0010002f60880000fffd;
mem[4382] = 80'h0010d8f0c0550102c000;
mem[4383] = 80'h00100001ffabffabffab;
mem[4384] = 80'h0010ff778b371e704403;
mem[4385] = 80'h0010e0afdbf5f5b6b66f;
mem[4386] = 80'h001068ad9463ace2603d;
mem[4387] = 80'h0111d000000000000000;
mem[4388] = 80'h00000000000000000000;
mem[4389] = 80'h10100000010000010010;
mem[4390] = 80'h00109400000208004500;
mem[4391] = 80'h0010002f60890000fffd;
mem[4392] = 80'h0010d8efc0550102c000;
mem[4393] = 80'h00100001ffabffabffab;
mem[4394] = 80'h0010ff76fae932a83dc1;
mem[4395] = 80'h00105f6409721843662e;
mem[4396] = 80'h001039e2a30bd0f422cd;
mem[4397] = 80'h0111a800000000000000;
mem[4398] = 80'h00000000000000000000;
mem[4399] = 80'h00000000000000000000;
mem[4400] = 80'h00000000000000000000;
mem[4401] = 80'h10100000010000010010;
mem[4402] = 80'h00109400000208004500;
mem[4403] = 80'h0010002f608a0000fffd;
mem[4404] = 80'h0010d8eec0550102c000;
mem[4405] = 80'h00100001ffabffabffab;
mem[4406] = 80'h0010ff75688b47c0b786;
mem[4407] = 80'h00109f387efa2e5d169d;
mem[4408] = 80'h0010cb2b825ee776925d;
mem[4409] = 80'h01115f00000000000000;
mem[4410] = 80'h00000000000000000000;
mem[4411] = 80'h00000000000000000000;
mem[4412] = 80'h00000000000000000000;
mem[4413] = 80'h10100000010000010010;
mem[4414] = 80'h00109400000208004500;
mem[4415] = 80'h0010002f608b0000fffd;
mem[4416] = 80'h0010d8edc0550102c000;
mem[4417] = 80'h00100001ffabffabffab;
mem[4418] = 80'h0010ff7419556b18ce44;
mem[4419] = 80'h001020f3ac7dc3a8c69d;
mem[4420] = 80'h00109a5a48c7727d6781;
mem[4421] = 80'h01113300000000000000;
mem[4422] = 80'h10100000010000010010;
mem[4423] = 80'h00109400000208004500;
mem[4424] = 80'h0010002f608c0000fffd;
mem[4425] = 80'h0010d8ecc0550102c000;
mem[4426] = 80'h00100001ffabffabffab;
mem[4427] = 80'h0010ff733d9181c9dacb;
mem[4428] = 80'h0010a04b436caf9427ee;
mem[4429] = 80'h00107f421de90d150407;
mem[4430] = 80'h0111a600000000000000;
mem[4431] = 80'h00000000000000000000;
mem[4432] = 80'h00000000000000000000;
mem[4433] = 80'h00000000000000000000;
mem[4434] = 80'h10100000010000010010;
mem[4435] = 80'h00109400000208004500;
mem[4436] = 80'h0010002f608d0000fffd;
mem[4437] = 80'h0010d8ebc0550102c000;
mem[4438] = 80'h00100001ffabffabffab;
mem[4439] = 80'h0010ff724c4fad11a309;
mem[4440] = 80'h00101f8091eb4261f76f;
mem[4441] = 80'h00102e1b7ecacbb6c900;
mem[4442] = 80'h01117800000000000000;
mem[4443] = 80'h00000000000000000000;
mem[4444] = 80'h10100000010000010010;
mem[4445] = 80'h00109400000208004500;
mem[4446] = 80'h0010002f608e0000fffd;
mem[4447] = 80'h0010d8eac0550102c000;
mem[4448] = 80'h00100001ffabffabffab;
mem[4449] = 80'h0010ff71de2dd879294e;
mem[4450] = 80'h0010dfdce663747f87fc;
mem[4451] = 80'h0010dcd4b906c7bb57b0;
mem[4452] = 80'h01111100000000000000;
mem[4453] = 80'h00000000000000000000;
mem[4454] = 80'h00000000000000000000;
mem[4455] = 80'h00000000000000000000;
mem[4456] = 80'h10100000010000010010;
mem[4457] = 80'h00109400000208004500;
mem[4458] = 80'h0010002f608f0000fffd;
mem[4459] = 80'h0010d8e9c0550102c000;
mem[4460] = 80'h00100001ffabffabffab;
mem[4461] = 80'h0010ff70aff3f4a1508c;
mem[4462] = 80'h0010601734e4998a57fd;
mem[4463] = 80'h00108d964253b4f27621;
mem[4464] = 80'h01115f00000000000000;
mem[4465] = 80'h00000000000000000000;
mem[4466] = 80'h10100000010000010010;
mem[4467] = 80'h00109400000208004500;
mem[4468] = 80'h0010002f60900000fffd;
mem[4469] = 80'h0010d8e8c0550102c000;
mem[4470] = 80'h00100001ffabffabffab;
mem[4471] = 80'h0010ff6fae822a8d88f5;
mem[4472] = 80'h0010a2a8ff291f67a201;
mem[4473] = 80'h0010e815cc3986eb8eeb;
mem[4474] = 80'h01111900000000000000;
mem[4475] = 80'h00000000000000000000;
mem[4476] = 80'h00000000000000000000;
mem[4477] = 80'h00000000000000000000;
mem[4478] = 80'h00000000000000000000;
mem[4479] = 80'h10100000010000010010;
mem[4480] = 80'h00109400000208004500;
mem[4481] = 80'h0010002f60910000fffd;
mem[4482] = 80'h0010d8e7c0550102c000;
mem[4483] = 80'h00100001ffabffabffab;
mem[4484] = 80'h0010ff6edf5c0655f137;
mem[4485] = 80'h00101d632daef2927383;
mem[4486] = 80'h0010b92ecc50f2a2b4e8;
mem[4487] = 80'h01116300000000000000;
mem[4488] = 80'h10100000010000010010;
mem[4489] = 80'h00109400000208004500;
mem[4490] = 80'h0010002f60920000fffd;
mem[4491] = 80'h0010d8e6c0550102c000;
mem[4492] = 80'h00100001ffabffabffab;
mem[4493] = 80'h0010ff6d4d3e733d7b70;
mem[4494] = 80'h0010dd3f5a26c48c0330;
mem[4495] = 80'h00104be7ed9b8b23cfde;
mem[4496] = 80'h0111ea00000000000000;
mem[4497] = 80'h00000000000000000000;
mem[4498] = 80'h00000000000000000000;
mem[4499] = 80'h00000000000000000000;
mem[4500] = 80'h10100000010000010010;
mem[4501] = 80'h00109400000208004500;
mem[4502] = 80'h0010002f60930000fffd;
mem[4503] = 80'h0010d8e5c0550102c000;
mem[4504] = 80'h00100001ffabffabffab;
mem[4505] = 80'h0010ff6c3ce05fe502b2;
mem[4506] = 80'h001062f488a12979d371;
mem[4507] = 80'h00101aa8daf28222b2eb;
mem[4508] = 80'h01110200000000000000;
mem[4509] = 80'h00000000000000000000;
mem[4510] = 80'h10100000010000010010;
mem[4511] = 80'h00109400000208004500;
mem[4512] = 80'h0010002f60940000fffd;
mem[4513] = 80'h0010d8e4c0550102c000;
mem[4514] = 80'h00100001ffabffabffab;
mem[4515] = 80'h0010ff6b1824b534163d;
mem[4516] = 80'h0010e24c67b045453242;
mem[4517] = 80'h0010ffbd43bc171e0cc8;
mem[4518] = 80'h0111d700000000000000;
mem[4519] = 80'h00000000000000000000;
mem[4520] = 80'h00000000000000000000;
mem[4521] = 80'h00000000000000000000;
mem[4522] = 80'h10100000010000010010;
mem[4523] = 80'h00109400000208004500;
mem[4524] = 80'h0010002f60950000fffd;
mem[4525] = 80'h0010d8e3c0550102c000;
mem[4526] = 80'h00100001ffabffabffab;
mem[4527] = 80'h0010ff6a69fa99ec6fff;
mem[4528] = 80'h00105d87b537a8b0e203;
mem[4529] = 80'h0010aef27448cb84fbfb;
mem[4530] = 80'h01113500000000000000;
mem[4531] = 80'h00000000000000000000;
mem[4532] = 80'h10100000010000010010;
mem[4533] = 80'h00109400000208004500;
mem[4534] = 80'h0010002f60960000fffd;
mem[4535] = 80'h0010d8e2c0550102c000;
mem[4536] = 80'h00100001ffabffabffab;
mem[4537] = 80'h0010ff69fb98ec84e5b8;
mem[4538] = 80'h00109ddbc2bf9eae9250;
mem[4539] = 80'h00105c2be7f95c65b828;
mem[4540] = 80'h0111ae00000000000000;
mem[4541] = 80'h00000000000000000000;
mem[4542] = 80'h00000000000000000000;
mem[4543] = 80'h00000000000000000000;
mem[4544] = 80'h00000000000000000000;
mem[4545] = 80'h10100000010000010010;
mem[4546] = 80'h00109400000208004500;
mem[4547] = 80'h0010002f60970000fffd;
mem[4548] = 80'h0010d8e1c0550102c000;
mem[4549] = 80'h00100001ffabffabffab;
mem[4550] = 80'h0010ff688a46c05c9c7a;
mem[4551] = 80'h001022101038735b4210;
mem[4552] = 80'h00100d57e16e42dd879a;
mem[4553] = 80'h01114300000000000000;
mem[4554] = 80'h10100000010000010010;
mem[4555] = 80'h00109400000208004500;
mem[4556] = 80'h0010002f60980000fffd;
mem[4557] = 80'h0010d8e0c0550102c000;
mem[4558] = 80'h00100001ffabffabffab;
mem[4559] = 80'h0010ff67b2113926cca7;
mem[4560] = 80'h00109caa1c9d46d750a6;
mem[4561] = 80'h0010973b2eb8318461fb;
mem[4562] = 80'h01118600000000000000;
mem[4563] = 80'h00000000000000000000;
mem[4564] = 80'h00000000000000000000;
mem[4565] = 80'h00000000000000000000;
mem[4566] = 80'h10100000010000010010;
mem[4567] = 80'h00109400000208004500;
mem[4568] = 80'h0010002f60990000fffd;
mem[4569] = 80'h0010d8dfc0550102c000;
mem[4570] = 80'h00100001ffabffabffab;
mem[4571] = 80'h0010ff66c3cf15feb565;
mem[4572] = 80'h00102361ce1aab2280e7;
mem[4573] = 80'h0010c674196b73b38ba8;
mem[4574] = 80'h01112100000000000000;
mem[4575] = 80'h00000000000000000000;
mem[4576] = 80'h10100000010000010010;
mem[4577] = 80'h00109400000208004500;
mem[4578] = 80'h0010002f609a0000fffd;
mem[4579] = 80'h0010d8dec0550102c000;
mem[4580] = 80'h00100001ffabffabffab;
mem[4581] = 80'h0010ff6551ad60963f22;
mem[4582] = 80'h0010e33db9929d3cf054;
mem[4583] = 80'h001034bd3815774ea798;
mem[4584] = 80'h01111f00000000000000;
mem[4585] = 80'h00000000000000000000;
mem[4586] = 80'h00000000000000000000;
mem[4587] = 80'h00000000000000000000;
mem[4588] = 80'h10100000010000010010;
mem[4589] = 80'h00109400000208004500;
mem[4590] = 80'h0010002f609b0000fffd;
mem[4591] = 80'h0010d8ddc0550102c000;
mem[4592] = 80'h00100001ffabffabffab;
mem[4593] = 80'h0010ff6420734c4e46e0;
mem[4594] = 80'h00105cf66b1570c927d5;
mem[4595] = 80'h00106561cbedba5137e2;
mem[4596] = 80'h0111ee00000000000000;
mem[4597] = 80'h00000000000000000000;
mem[4598] = 80'h00000000000000000000;
mem[4599] = 80'h00000000000000000000;
mem[4600] = 80'h10100000010000010010;
mem[4601] = 80'h00109400000208004500;
mem[4602] = 80'h0010002f609c0000fffd;
mem[4603] = 80'h0010d8dcc0550102c000;
mem[4604] = 80'h00100001ffabffabffab;
mem[4605] = 80'h0010ff6304b7a69f526f;
mem[4606] = 80'h0010dc4e84041cf5c6a6;
mem[4607] = 80'h001080799e6d9fb47d5e;
mem[4608] = 80'h0111c000000000000000;
mem[4609] = 80'h00000000000000000000;
mem[4610] = 80'h10100000010000010010;
mem[4611] = 80'h00109400000208004500;
mem[4612] = 80'h0010002f609d0000fffd;
mem[4613] = 80'h0010d8dbc0550102c000;
mem[4614] = 80'h00100001ffabffabffab;
mem[4615] = 80'h0010ff6275698a472bad;
mem[4616] = 80'h001063855683f10016a0;
mem[4617] = 80'h0010d1a2f2f24e89c943;
mem[4618] = 80'h01119a00000000000000;
mem[4619] = 80'h00000000000000000000;
mem[4620] = 80'h10100000010000010010;
mem[4621] = 80'h00109400000208004500;
mem[4622] = 80'h0010002f609e0000fffd;
mem[4623] = 80'h0010d8dac0550102c000;
mem[4624] = 80'h00100001ffabffabffab;
mem[4625] = 80'h0010ff61e70bff2fa1ea;
mem[4626] = 80'h0010a3d9210bc71e662b;
mem[4627] = 80'h001023e7ef6172fc4076;
mem[4628] = 80'h01110500000000000000;
mem[4629] = 80'h00000000000000000000;
mem[4630] = 80'h00000000000000000000;
mem[4631] = 80'h00000000000000000000;
mem[4632] = 80'h00000000000000000000;
mem[4633] = 80'h10100000010000010010;
mem[4634] = 80'h00109400000208004500;
mem[4635] = 80'h0010002f609f0000fffd;
mem[4636] = 80'h0010d8d9c0550102c000;
mem[4637] = 80'h00100001ffabffabffab;
mem[4638] = 80'h0010ff6096d5d3f7d828;
mem[4639] = 80'h00101c12f38c2aebb6b2;
mem[4640] = 80'h00107234563803d4048b;
mem[4641] = 80'h01118e00000000000000;
mem[4642] = 80'h00000000000000000000;
mem[4643] = 80'h10100000010000010010;
mem[4644] = 80'h00109400000208004500;
mem[4645] = 80'h0010002f60a00000fffd;
mem[4646] = 80'h0010d8d8c0550102c000;
mem[4647] = 80'h00100001ffabffabffab;
mem[4648] = 80'h0010ff5fe5e843761119;
mem[4649] = 80'h001026a6b690cac58d53;
mem[4650] = 80'h0010e9eb4aec5bda9454;
mem[4651] = 80'h01118c00000000000000;
mem[4652] = 80'h00000000000000000000;
mem[4653] = 80'h00000000000000000000;
mem[4654] = 80'h00000000000000000000;
mem[4655] = 80'h10100000010000010010;
mem[4656] = 80'h00109400000208004500;
mem[4657] = 80'h0010002f60a10000fffd;
mem[4658] = 80'h0010d8d7c0550102c000;
mem[4659] = 80'h00100001ffabffabffab;
mem[4660] = 80'h0010ff5e94366fae68db;
mem[4661] = 80'h0010996d641727305d5a;
mem[4662] = 80'h0010b82018b1407b222e;
mem[4663] = 80'h0111ab00000000000000;
mem[4664] = 80'h00000000000000000000;
mem[4665] = 80'h10100000010000010010;
mem[4666] = 80'h00109400000208004500;
mem[4667] = 80'h0010002f60a20000fffd;
mem[4668] = 80'h0010d8d6c0550102c000;
mem[4669] = 80'h00100001ffabffabffab;
mem[4670] = 80'h0010ff5d06541ac6e29c;
mem[4671] = 80'h00105931139f112e2dd1;
mem[4672] = 80'h00104a6505b70046e89e;
mem[4673] = 80'h01116100000000000000;
mem[4674] = 80'h00000000000000000000;
mem[4675] = 80'h00000000000000000000;
mem[4676] = 80'h00000000000000000000;
mem[4677] = 80'h10100000010000010010;
mem[4678] = 80'h00109400000208004500;
mem[4679] = 80'h0010002f60a30000fffd;
mem[4680] = 80'h0010d8d5c0550102c000;
mem[4681] = 80'h00100001ffabffabffab;
mem[4682] = 80'h0010ff5c778a361e9b5e;
mem[4683] = 80'h0010e6fac118fcdbfda8;
mem[4684] = 80'h00101ba60e5deaba7dd1;
mem[4685] = 80'h0111c200000000000000;
mem[4686] = 80'h00000000000000000000;
mem[4687] = 80'h10100000010000010010;
mem[4688] = 80'h00109400000208004500;
mem[4689] = 80'h0010002f60a40000fffd;
mem[4690] = 80'h0010d8d4c0550102c000;
mem[4691] = 80'h00100001ffabffabffab;
mem[4692] = 80'h0010ff5b534edccf8fd1;
mem[4693] = 80'h001066422e0990e71d12;
mem[4694] = 80'h0010fe25a749587fd624;
mem[4695] = 80'h0111d100000000000000;
mem[4696] = 80'h00000000000000000000;
mem[4697] = 80'h00000000000000000000;
mem[4698] = 80'h00000000000000000000;
mem[4699] = 80'h10100000010000010010;
mem[4700] = 80'h00109400000208004500;
mem[4701] = 80'h0010002f60a50000fffd;
mem[4702] = 80'h0010d8d3c0550102c000;
mem[4703] = 80'h00100001ffabffabffab;
mem[4704] = 80'h0010ff5a2290f017f613;
mem[4705] = 80'h0010d989fc8e7d12cd5b;
mem[4706] = 80'h0010afe3397eeda76105;
mem[4707] = 80'h01114d00000000000000;
mem[4708] = 80'h00000000000000000000;
mem[4709] = 80'h10100000010000010010;
mem[4710] = 80'h00109400000208004500;
mem[4711] = 80'h0010002f60a60000fffd;
mem[4712] = 80'h0010d8d2c0550102c000;
mem[4713] = 80'h00100001ffabffabffab;
mem[4714] = 80'h0010ff59b0f2857f7c54;
mem[4715] = 80'h001019d58b064b0cbd90;
mem[4716] = 80'h00105dabe8bb5987a435;
mem[4717] = 80'h0111b800000000000000;
mem[4718] = 80'h00000000000000000000;
mem[4719] = 80'h00000000000000000000;
mem[4720] = 80'h00000000000000000000;
mem[4721] = 80'h10100000010000010010;
mem[4722] = 80'h00109400000208004500;
mem[4723] = 80'h0010002f60a70000fffd;
mem[4724] = 80'h0010d8d1c0550102c000;
mem[4725] = 80'h00100001ffabffabffab;
mem[4726] = 80'h0010ff58c12ca9a70596;
mem[4727] = 80'h0010a61e5981a6f96dc9;
mem[4728] = 80'h00100c6e056c69f7b43c;
mem[4729] = 80'h01119800000000000000;
mem[4730] = 80'h00000000000000000000;
mem[4731] = 80'h10100000010000010010;
mem[4732] = 80'h00109400000208004500;
mem[4733] = 80'h0010002f60a80000fffd;
mem[4734] = 80'h0010d8d0c0550102c000;
mem[4735] = 80'h00100001ffabffabffab;
mem[4736] = 80'h0010ff57f97b50dd554b;
mem[4737] = 80'h001018a4552493757ff7;
mem[4738] = 80'h00109690fb3d4d48a893;
mem[4739] = 80'h01111c00000000000000;
mem[4740] = 80'h00000000000000000000;
mem[4741] = 80'h10100000010000010010;
mem[4742] = 80'h00109400000208004500;
mem[4743] = 80'h0010002f60a90000fffd;
mem[4744] = 80'h0010d8cfc0550102c000;
mem[4745] = 80'h00100001ffabffabffab;
mem[4746] = 80'h0010ff5688a57c052c89;
mem[4747] = 80'h0010a76f87a37e80afbe;
mem[4748] = 80'h0010c75665cc448d4324;
mem[4749] = 80'h01114e00000000000000;
mem[4750] = 80'h00000000000000000000;
mem[4751] = 80'h00000000000000000000;
mem[4752] = 80'h00000000000000000000;
mem[4753] = 80'h10100000010000010010;
mem[4754] = 80'h00109400000208004500;
mem[4755] = 80'h0010002f60aa0000fffd;
mem[4756] = 80'h0010d8cec0550102c000;
mem[4757] = 80'h00100001ffabffabffab;
mem[4758] = 80'h0010ff551ac7096da6ce;
mem[4759] = 80'h00106733f02b489edf76;
mem[4760] = 80'h0010354be7e79872ac3d;
mem[4761] = 80'h01112c00000000000000;
mem[4762] = 80'h00000000000000000000;
mem[4763] = 80'h00000000000000000000;
mem[4764] = 80'h00000000000000000000;
mem[4765] = 80'h10100000010000010010;
mem[4766] = 80'h00109400000208004500;
mem[4767] = 80'h0010002f60ab0000fffd;
mem[4768] = 80'h0010d8cdc0550102c000;
mem[4769] = 80'h00100001ffabffabffab;
mem[4770] = 80'h0010ff546b1925b5df0c;
mem[4771] = 80'h0010d8f822aca56b0f0f;
mem[4772] = 80'h00106488ec278f077b15;
mem[4773] = 80'h01112300000000000000;
mem[4774] = 80'h10100000010000010010;
mem[4775] = 80'h00109400000208004500;
mem[4776] = 80'h0010002f60ac0000fffd;
mem[4777] = 80'h0010d8ccc0550102c000;
mem[4778] = 80'h00100001ffabffabffab;
mem[4779] = 80'h0010ff534fddcf64cb83;
mem[4780] = 80'h00105840cdbdc957ee74;
mem[4781] = 80'h001081191002a65628c4;
mem[4782] = 80'h01117d00000000000000;
mem[4783] = 80'h00000000000000000000;
mem[4784] = 80'h00000000000000000000;
mem[4785] = 80'h00000000000000000000;
mem[4786] = 80'h10100000010000010010;
mem[4787] = 80'h00109400000208004500;
mem[4788] = 80'h0010002f60ad0000fffd;
mem[4789] = 80'h0010d8cbc0550102c000;
mem[4790] = 80'h00100001ffabffabffab;
mem[4791] = 80'h0010ff523e03e3bcb241;
mem[4792] = 80'h0010e78b1f3a24a23dfd;
mem[4793] = 80'h0010d0908ab5677e5670;
mem[4794] = 80'h01116900000000000000;
mem[4795] = 80'h00000000000000000000;
mem[4796] = 80'h10100000010000010010;
mem[4797] = 80'h00109400000208004500;
mem[4798] = 80'h0010002f60ae0000fffd;
mem[4799] = 80'h0010d8cac0550102c000;
mem[4800] = 80'h00100001ffabffabffab;
mem[4801] = 80'h0010ff51ac6196d43806;
mem[4802] = 80'h001027d768b212bc4d76;
mem[4803] = 80'h001022d597e0d9cf4d53;
mem[4804] = 80'h01116800000000000000;
mem[4805] = 80'h00000000000000000000;
mem[4806] = 80'h00000000000000000000;
mem[4807] = 80'h00000000000000000000;
mem[4808] = 80'h10100000010000010010;
mem[4809] = 80'h00109400000208004500;
mem[4810] = 80'h0010002f60af0000fffd;
mem[4811] = 80'h0010d8c9c0550102c000;
mem[4812] = 80'h00100001ffabffabffab;
mem[4813] = 80'h0010ff50ddbfba0c41c4;
mem[4814] = 80'h0010981cba35ff499d6f;
mem[4815] = 80'h0010731db6f50d877376;
mem[4816] = 80'h01117300000000000000;
mem[4817] = 80'h00000000000000000000;
mem[4818] = 80'h10100000010000010010;
mem[4819] = 80'h00109400000208004500;
mem[4820] = 80'h0010002f60b00000fffd;
mem[4821] = 80'h0010d8c8c0550102c000;
mem[4822] = 80'h00100001ffabffabffab;
mem[4823] = 80'h0010ff4fdcce642099bd;
mem[4824] = 80'h00105aa371f879a4689a;
mem[4825] = 80'h00101624a004c0bc21cb;
mem[4826] = 80'h01112c00000000000000;
mem[4827] = 80'h00000000000000000000;
mem[4828] = 80'h00000000000000000000;
mem[4829] = 80'h00000000000000000000;
mem[4830] = 80'h00000000000000000000;
mem[4831] = 80'h10100000010000010010;
mem[4832] = 80'h00109400000208004500;
mem[4833] = 80'h0010002f60b10000fffd;
mem[4834] = 80'h0010d8c7c0550102c000;
mem[4835] = 80'h00100001ffabffabffab;
mem[4836] = 80'h0010ff4ead1048f8e07f;
mem[4837] = 80'h0010e568a37f9451b813;
mem[4838] = 80'h001047f46ae6a1469094;
mem[4839] = 80'h0111b200000000000000;
mem[4840] = 80'h10100000010000010010;
mem[4841] = 80'h00109400000208004500;
mem[4842] = 80'h0010002f60b20000fffd;
mem[4843] = 80'h0010d8c6c0550102c000;
mem[4844] = 80'h00100001ffabffabffab;
mem[4845] = 80'h0010ff4d3f723d906a38;
mem[4846] = 80'h00102534d4f7a24fc898;
mem[4847] = 80'h0010b5b177b18695c252;
mem[4848] = 80'h01110800000000000000;
mem[4849] = 80'h00000000000000000000;
mem[4850] = 80'h00000000000000000000;
mem[4851] = 80'h00000000000000000000;
mem[4852] = 80'h10100000010000010010;
mem[4853] = 80'h00109400000208004500;
mem[4854] = 80'h0010002f60b30000fffd;
mem[4855] = 80'h0010d8c5c0550102c000;
mem[4856] = 80'h00100001ffabffabffab;
mem[4857] = 80'h0010ff4c4eac114813fa;
mem[4858] = 80'h00109aff06704fba18e1;
mem[4859] = 80'h0010e4727c4721193707;
mem[4860] = 80'h01114500000000000000;
mem[4861] = 80'h00000000000000000000;
mem[4862] = 80'h10100000010000010010;
mem[4863] = 80'h00109400000208004500;
mem[4864] = 80'h0010002f60b40000fffd;
mem[4865] = 80'h0010d8c4c0550102c000;
mem[4866] = 80'h00100001ffabffabffab;
mem[4867] = 80'h0010ff4b6a68fb990775;
mem[4868] = 80'h00101a47e9612386f9da;
mem[4869] = 80'h001001ee4c4523f89228;
mem[4870] = 80'h01110800000000000000;
mem[4871] = 80'h00000000000000000000;
mem[4872] = 80'h00000000000000000000;
mem[4873] = 80'h00000000000000000000;
mem[4874] = 80'h10100000010000010010;
mem[4875] = 80'h00109400000208004500;
mem[4876] = 80'h0010002f60b50000fffd;
mem[4877] = 80'h0010d8c3c0550102c000;
mem[4878] = 80'h00100001ffabffabffab;
mem[4879] = 80'h0010ff4a1bb6d7417eb7;
mem[4880] = 80'h0010a58c3be6ce732993;
mem[4881] = 80'h00105028d2639229c2bd;
mem[4882] = 80'h0111c000000000000000;
mem[4883] = 80'h00000000000000000000;
mem[4884] = 80'h10100000010000010010;
mem[4885] = 80'h00109400000208004500;
mem[4886] = 80'h0010002f60b60000fffd;
mem[4887] = 80'h0010d8c2c0550102c000;
mem[4888] = 80'h00100001ffabffabffab;
mem[4889] = 80'h0010ff4989d4a229f4f0;
mem[4890] = 80'h001065d04c6ef86d58df;
mem[4891] = 80'h0010a2d53c65fc9f8b05;
mem[4892] = 80'h01111300000000000000;
mem[4893] = 80'h00000000000000000000;
mem[4894] = 80'h00000000000000000000;
mem[4895] = 80'h00000000000000000000;
mem[4896] = 80'h00000000000000000000;
mem[4897] = 80'h10100000010000010010;
mem[4898] = 80'h00109400000208004500;
mem[4899] = 80'h0010002f60b70000fffd;
mem[4900] = 80'h0010d8c1c0550102c000;
mem[4901] = 80'h00100001ffabffabffab;
mem[4902] = 80'h0010ff48f80a8ef18d32;
mem[4903] = 80'h0010da1b9ee91598889e;
mem[4904] = 80'h0010f39a0bb1d5a30635;
mem[4905] = 80'h01119100000000000000;
mem[4906] = 80'h10100000010000010010;
mem[4907] = 80'h00109400000208004500;
mem[4908] = 80'h0010002f60b80000fffd;
mem[4909] = 80'h0010d8c0c0550102c000;
mem[4910] = 80'h00100001ffabffabffab;
mem[4911] = 80'h0010ff47c05d778bddef;
mem[4912] = 80'h001064a1924c20149a38;
mem[4913] = 80'h001069f5b7af17da45c5;
mem[4914] = 80'h0111ac00000000000000;
mem[4915] = 80'h00000000000000000000;
mem[4916] = 80'h00000000000000000000;
mem[4917] = 80'h00000000000000000000;
mem[4918] = 80'h10100000010000010010;
mem[4919] = 80'h00109400000208004500;
mem[4920] = 80'h0010002f60b90000fffd;
mem[4921] = 80'h0010d8bfc0550102c000;
mem[4922] = 80'h00100001ffabffabffab;
mem[4923] = 80'h0010ff46b1835b53a42d;
mem[4924] = 80'h0010db6a40cbcde14a79;
mem[4925] = 80'h001038ba806961be3870;
mem[4926] = 80'h01112e00000000000000;
mem[4927] = 80'h00000000000000000000;
mem[4928] = 80'h10100000010000010010;
mem[4929] = 80'h00109400000208004500;
mem[4930] = 80'h0010002f60ba0000fffd;
mem[4931] = 80'h0010d8bec0550102c000;
mem[4932] = 80'h00100001ffabffabffab;
mem[4933] = 80'h0010ff4523e12e3b2e6a;
mem[4934] = 80'h00101b363743fbff3a3a;
mem[4935] = 80'h0010ca60601fcc1898c0;
mem[4936] = 80'h0111b000000000000000;
mem[4937] = 80'h00000000000000000000;
mem[4938] = 80'h00000000000000000000;
mem[4939] = 80'h00000000000000000000;
mem[4940] = 80'h10100000010000010010;
mem[4941] = 80'h00109400000208004500;
mem[4942] = 80'h0010002f60bb0000fffd;
mem[4943] = 80'h0010d8bdc0550102c000;
mem[4944] = 80'h00100001ffabffabffab;
mem[4945] = 80'h0010ff44523f02e357a8;
mem[4946] = 80'h0010a4fde5c4160aea7b;
mem[4947] = 80'h00109b2f5778d5f3d8c1;
mem[4948] = 80'h0111db00000000000000;
mem[4949] = 80'h00000000000000000000;
mem[4950] = 80'h00000000000000000000;
mem[4951] = 80'h00000000000000000000;
mem[4952] = 80'h10100000010000010010;
mem[4953] = 80'h00109400000208004500;
mem[4954] = 80'h0010002f60bc0000fffd;
mem[4955] = 80'h0010d8bcc0550102c000;
mem[4956] = 80'h00100001ffabffabffab;
mem[4957] = 80'h0010ff4376fbe8324327;
mem[4958] = 80'h001024450ad57a360b38;
mem[4959] = 80'h00107e3297ab93e7212c;
mem[4960] = 80'h01117800000000000000;
mem[4961] = 80'h00000000000000000000;
mem[4962] = 80'h10100000010000010010;
mem[4963] = 80'h00109400000208004500;
mem[4964] = 80'h0010002f60bd0000fffd;
mem[4965] = 80'h0010d8bbc0550102c000;
mem[4966] = 80'h00100001ffabffabffab;
mem[4967] = 80'h0010ff420725c4ea3ae5;
mem[4968] = 80'h00109b8ed85297c3db38;
mem[4969] = 80'h00102f435da785be2027;
mem[4970] = 80'h01115400000000000000;
mem[4971] = 80'h00000000000000000000;
mem[4972] = 80'h10100000010000010010;
mem[4973] = 80'h00109400000208004500;
mem[4974] = 80'h0010002f60be0000fffd;
mem[4975] = 80'h0010d8bac0550102c000;
mem[4976] = 80'h00100001ffabffabffab;
mem[4977] = 80'h0010ff419547b182b0a2;
mem[4978] = 80'h00105bd2afdaa1ddabbb;
mem[4979] = 80'h0010dd8fe97ae811b72f;
mem[4980] = 80'h01111300000000000000;
mem[4981] = 80'h00000000000000000000;
mem[4982] = 80'h00000000000000000000;
mem[4983] = 80'h00000000000000000000;
mem[4984] = 80'h00000000000000000000;
mem[4985] = 80'h10100000010000010010;
mem[4986] = 80'h00109400000208004500;
mem[4987] = 80'h0010002f60bf0000fffd;
mem[4988] = 80'h0010d8b9c0550102c000;
mem[4989] = 80'h00100001ffabffabffab;
mem[4990] = 80'h0010ff40e4999d5ac960;
mem[4991] = 80'h0010e4197d5d4c28743a;
mem[4992] = 80'h00108cfabb954aeef0ed;
mem[4993] = 80'h0111e100000000000000;
mem[4994] = 80'h00000000000000000000;
mem[4995] = 80'h10100000010000010010;
mem[4996] = 80'h00109400000208004500;
mem[4997] = 80'h0010002f60c00000fffd;
mem[4998] = 80'h0010d8b8c0550102c000;
mem[4999] = 80'h00100001ffabffabffab;
mem[5000] = 80'h0010ff3f733c908122c0;
mem[5001] = 80'h00102eba25e36181d3e8;
mem[5002] = 80'h0010eb152a253a4dc47c;
mem[5003] = 80'h01117e00000000000000;
mem[5004] = 80'h00000000000000000000;
mem[5005] = 80'h00000000000000000000;
mem[5006] = 80'h00000000000000000000;
mem[5007] = 80'h10100000010000010010;
mem[5008] = 80'h00109400000208004500;
mem[5009] = 80'h0010002f60c10000fffd;
mem[5010] = 80'h0010d8b7c0550102c000;
mem[5011] = 80'h00100001ffabffabffab;
mem[5012] = 80'h0010ff3e02e2bc595b02;
mem[5013] = 80'h00109171f7648c7403e9;
mem[5014] = 80'h0010ba57d1f74095ba03;
mem[5015] = 80'h01117500000000000000;
mem[5016] = 80'h00000000000000000000;
mem[5017] = 80'h10100000010000010010;
mem[5018] = 80'h00109400000208004500;
mem[5019] = 80'h0010002f60c20000fffd;
mem[5020] = 80'h0010d8b6c0550102c000;
mem[5021] = 80'h00100001ffabffabffab;
mem[5022] = 80'h0010ff3d9080c931d145;
mem[5023] = 80'h0010512d80ecba6a736a;
mem[5024] = 80'h0010489b6540270947cc;
mem[5025] = 80'h01114d00000000000000;
mem[5026] = 80'h00000000000000000000;
mem[5027] = 80'h00000000000000000000;
mem[5028] = 80'h00000000000000000000;
mem[5029] = 80'h10100000010000010010;
mem[5030] = 80'h00109400000208004500;
mem[5031] = 80'h0010002f60c30000fffd;
mem[5032] = 80'h0010d8b5c0550102c000;
mem[5033] = 80'h00100001ffabffabffab;
mem[5034] = 80'h0010ff3ce15ee5e9a887;
mem[5035] = 80'h0010eee6526b579fa3e8;
mem[5036] = 80'h001019975581e40baa04;
mem[5037] = 80'h0111a300000000000000;
mem[5038] = 80'h00000000000000000000;
mem[5039] = 80'h10100000010000010010;
mem[5040] = 80'h00109400000208004500;
mem[5041] = 80'h0010002f60c40000fffd;
mem[5042] = 80'h0010d8b4c0550102c000;
mem[5043] = 80'h00100001ffabffabffab;
mem[5044] = 80'h0010ff3bc59a0f38bc08;
mem[5045] = 80'h00106e5ebd7a3ba342ab;
mem[5046] = 80'h0010fc8a9536336e5e70;
mem[5047] = 80'h01118600000000000000;
mem[5048] = 80'h00000000000000000000;
mem[5049] = 80'h00000000000000000000;
mem[5050] = 80'h00000000000000000000;
mem[5051] = 80'h10100000010000010010;
mem[5052] = 80'h00109400000208004500;
mem[5053] = 80'h0010002f60c50000fffd;
mem[5054] = 80'h0010d8b3c0550102c000;
mem[5055] = 80'h00100001ffabffabffab;
mem[5056] = 80'h0010ff3ab44423e0c5ca;
mem[5057] = 80'h0010d1956ffdd65692ea;
mem[5058] = 80'h0010adc5a23b6712f85e;
mem[5059] = 80'h01114200000000000000;
mem[5060] = 80'h00000000000000000000;
mem[5061] = 80'h10100000010000010010;
mem[5062] = 80'h00109400000208004500;
mem[5063] = 80'h0010002f60c60000fffd;
mem[5064] = 80'h0010d8b2c0550102c000;
mem[5065] = 80'h00100001ffabffabffab;
mem[5066] = 80'h0010ff39262656884f8d;
mem[5067] = 80'h001011c91875e048e229;
mem[5068] = 80'h00105f04dad50dbb22de;
mem[5069] = 80'h01110a00000000000000;
mem[5070] = 80'h00000000000000000000;
mem[5071] = 80'h00000000000000000000;
mem[5072] = 80'h00000000000000000000;
mem[5073] = 80'h10100000010000010010;
mem[5074] = 80'h00109400000208004500;
mem[5075] = 80'h0010002f60c70000fffd;
mem[5076] = 80'h0010d8b1c0550102c000;
mem[5077] = 80'h00100001ffabffabffab;
mem[5078] = 80'h0010ff3857f87a50364f;
mem[5079] = 80'h0010ae02caf20dbd3268;
mem[5080] = 80'h00100e4bedc942ac361c;
mem[5081] = 80'h01112f00000000000000;
mem[5082] = 80'h00000000000000000000;
mem[5083] = 80'h10100000010000010010;
mem[5084] = 80'h00109400000208004500;
mem[5085] = 80'h0010002f60c80000fffd;
mem[5086] = 80'h0010d8b0c0550102c000;
mem[5087] = 80'h00100001ffabffabffab;
mem[5088] = 80'h0010ff376faf832a6692;
mem[5089] = 80'h001010b8c6573831214e;
mem[5090] = 80'h00109408f9c3e8d84863;
mem[5091] = 80'h0111fa00000000000000;
mem[5092] = 80'h00000000000000000000;
mem[5093] = 80'h10100000010000010010;
mem[5094] = 80'h00109400000208004500;
mem[5095] = 80'h0010002f60c90000fffd;
mem[5096] = 80'h0010d8afc0550102c000;
mem[5097] = 80'h00100001ffabffabffab;
mem[5098] = 80'h0010ff361e71aff21f50;
mem[5099] = 80'h0010af7314d0d5c4f10e;
mem[5100] = 80'h0010c574ff88c2238259;
mem[5101] = 80'h0111b200000000000000;
mem[5102] = 80'h00000000000000000000;
mem[5103] = 80'h00000000000000000000;
mem[5104] = 80'h00000000000000000000;
mem[5105] = 80'h10100000010000010010;
mem[5106] = 80'h00109400000208004500;
mem[5107] = 80'h0010002f60ca0000fffd;
mem[5108] = 80'h0010d8aec0550102c000;
mem[5109] = 80'h00100001ffabffabffab;
mem[5110] = 80'h0010ff358c13da9a9517;
mem[5111] = 80'h00106f2f6358e3da81cd;
mem[5112] = 80'h001037b5871f0d52cd98;
mem[5113] = 80'h0111a200000000000000;
mem[5114] = 80'h00000000000000000000;
mem[5115] = 80'h00000000000000000000;
mem[5116] = 80'h00000000000000000000;
mem[5117] = 80'h10100000010000010010;
mem[5118] = 80'h00109400000208004500;
mem[5119] = 80'h0010002f60cb0000fffd;
mem[5120] = 80'h0010d8adc0550102c000;
mem[5121] = 80'h00100001ffabffabffab;
mem[5122] = 80'h0010ff34fdcdf642ecd5;
mem[5123] = 80'h0010d0e4b1df0e2f518c;
mem[5124] = 80'h001066fab06a2550fdb3;
mem[5125] = 80'h0111e000000000000000;
mem[5126] = 80'h10100000010000010010;
mem[5127] = 80'h00109400000208004500;
mem[5128] = 80'h0010002f60cc0000fffd;
mem[5129] = 80'h0010d8acc0550102c000;
mem[5130] = 80'h00100001ffabffabffab;
mem[5131] = 80'h0010ff33d9091c93f85a;
mem[5132] = 80'h0010505c5ece6213b0cf;
mem[5133] = 80'h001083e770df5bfb70fb;
mem[5134] = 80'h01115800000000000000;
mem[5135] = 80'h00000000000000000000;
mem[5136] = 80'h00000000000000000000;
mem[5137] = 80'h00000000000000000000;
mem[5138] = 80'h10100000010000010010;
mem[5139] = 80'h00109400000208004500;
mem[5140] = 80'h0010002f60cd0000fffd;
mem[5141] = 80'h0010d8abc0550102c000;
mem[5142] = 80'h00100001ffabffabffab;
mem[5143] = 80'h0010ff32a8d7304b8198;
mem[5144] = 80'h0010ef978c498fe6604e;
mem[5145] = 80'h0010d2be133d53e0b4c1;
mem[5146] = 80'h01112800000000000000;
mem[5147] = 80'h00000000000000000000;
mem[5148] = 80'h10100000010000010010;
mem[5149] = 80'h00109400000208004500;
mem[5150] = 80'h0010002f60ce0000fffd;
mem[5151] = 80'h0010d8aac0550102c000;
mem[5152] = 80'h00100001ffabffabffab;
mem[5153] = 80'h0010ff313ab545230bdf;
mem[5154] = 80'h00102fcbfbc1b9f810cd;
mem[5155] = 80'h00102072a751b6a4b774;
mem[5156] = 80'h01117100000000000000;
mem[5157] = 80'h00000000000000000000;
mem[5158] = 80'h00000000000000000000;
mem[5159] = 80'h00000000000000000000;
mem[5160] = 80'h10100000010000010010;
mem[5161] = 80'h00109400000208004500;
mem[5162] = 80'h0010002f60cf0000fffd;
mem[5163] = 80'h0010d8a9c0550102c000;
mem[5164] = 80'h00100001ffabffabffab;
mem[5165] = 80'h0010ff304b6b69fb721d;
mem[5166] = 80'h001090002946540dc0cb;
mem[5167] = 80'h001071a9cb81cd3242db;
mem[5168] = 80'h01115200000000000000;
mem[5169] = 80'h00000000000000000000;
mem[5170] = 80'h10100000010000010010;
mem[5171] = 80'h00109400000208004500;
mem[5172] = 80'h0010002f60d00000fffd;
mem[5173] = 80'h0010d8a8c0550102c000;
mem[5174] = 80'h00100001ffabffabffab;
mem[5175] = 80'h0010ff2f4a1ab7d7aa64;
mem[5176] = 80'h001052bfe28bd2e0353f;
mem[5177] = 80'h001014a3ec6b153534e6;
mem[5178] = 80'h0111c500000000000000;
mem[5179] = 80'h00000000000000000000;
mem[5180] = 80'h00000000000000000000;
mem[5181] = 80'h00000000000000000000;
mem[5182] = 80'h00000000000000000000;
mem[5183] = 80'h10100000010000010010;
mem[5184] = 80'h00109400000208004500;
mem[5185] = 80'h0010002f60d10000fffd;
mem[5186] = 80'h0010d8a7c0550102c000;
mem[5187] = 80'h00100001ffabffabffab;
mem[5188] = 80'h0010ff2e3bc49b0fd3a6;
mem[5189] = 80'h0010ed74300c3f15e6a6;
mem[5190] = 80'h0010452905f0c73faaa9;
mem[5191] = 80'h01115b00000000000000;
mem[5192] = 80'h10100000010000010010;
mem[5193] = 80'h00109400000208004500;
mem[5194] = 80'h0010002f60d20000fffd;
mem[5195] = 80'h0010d8a6c0550102c000;
mem[5196] = 80'h00100001ffabffabffab;
mem[5197] = 80'h0010ff2da9a6ee6759e1;
mem[5198] = 80'h00102d284784090b962d;
mem[5199] = 80'h0010b76c18912a3742c2;
mem[5200] = 80'h01111300000000000000;
mem[5201] = 80'h00000000000000000000;
mem[5202] = 80'h00000000000000000000;
mem[5203] = 80'h00000000000000000000;
mem[5204] = 80'h10100000010000010010;
mem[5205] = 80'h00109400000208004500;
mem[5206] = 80'h0010002f60d30000fffd;
mem[5207] = 80'h0010d8a5c0550102c000;
mem[5208] = 80'h00100001ffabffabffab;
mem[5209] = 80'h0010ff2cd878c2bf2023;
mem[5210] = 80'h001092e39503e4fe4624;
mem[5211] = 80'h0010e6a74ac5c0ec6430;
mem[5212] = 80'h01116700000000000000;
mem[5213] = 80'h00000000000000000000;
mem[5214] = 80'h10100000010000010010;
mem[5215] = 80'h00109400000208004500;
mem[5216] = 80'h0010002f60d40000fffd;
mem[5217] = 80'h0010d8a4c0550102c000;
mem[5218] = 80'h00100001ffabffabffab;
mem[5219] = 80'h0010ff2bfcbc286e34ac;
mem[5220] = 80'h0010125b7a1288c2a75f;
mem[5221] = 80'h00100336b63730150e97;
mem[5222] = 80'h01110800000000000000;
mem[5223] = 80'h00000000000000000000;
mem[5224] = 80'h00000000000000000000;
mem[5225] = 80'h00000000000000000000;
mem[5226] = 80'h10100000010000010010;
mem[5227] = 80'h00109400000208004500;
mem[5228] = 80'h0010002f60d50000fffd;
mem[5229] = 80'h0010d8a3c0550102c000;
mem[5230] = 80'h00100001ffabffabffab;
mem[5231] = 80'h0010ff2a8d6204b64d6e;
mem[5232] = 80'h0010ad90a89565377726;
mem[5233] = 80'h001052f5bdd4dd94ed2e;
mem[5234] = 80'h0111dc00000000000000;
mem[5235] = 80'h00000000000000000000;
mem[5236] = 80'h10100000010000010010;
mem[5237] = 80'h00109400000208004500;
mem[5238] = 80'h0010002f60d60000fffd;
mem[5239] = 80'h0010d8a2c0550102c000;
mem[5240] = 80'h00100001ffabffabffab;
mem[5241] = 80'h0010ff291f0071dec729;
mem[5242] = 80'h00106dccdf1d5329076c;
mem[5243] = 80'h0010a095c5b89af1aaac;
mem[5244] = 80'h01111400000000000000;
mem[5245] = 80'h00000000000000000000;
mem[5246] = 80'h00000000000000000000;
mem[5247] = 80'h00000000000000000000;
mem[5248] = 80'h00000000000000000000;
mem[5249] = 80'h10100000010000010010;
mem[5250] = 80'h00109400000208004500;
mem[5251] = 80'h0010002f60d70000fffd;
mem[5252] = 80'h0010d8a1c0550102c000;
mem[5253] = 80'h00100001ffabffabffab;
mem[5254] = 80'h0010ff286ede5d06beeb;
mem[5255] = 80'h0010d2070d9abedcd725;
mem[5256] = 80'h0010f1535b0eb3db33fc;
mem[5257] = 80'h01116b00000000000000;
mem[5258] = 80'h10100000010000010010;
mem[5259] = 80'h00109400000208004500;
mem[5260] = 80'h0010002f60d80000fffd;
mem[5261] = 80'h0010d8a0c0550102c000;
mem[5262] = 80'h00100001ffabffabffab;
mem[5263] = 80'h0010ff275689a47cee36;
mem[5264] = 80'h00106cbd013f8b50c59b;
mem[5265] = 80'h00106bb63dfcae4865d4;
mem[5266] = 80'h01115f00000000000000;
mem[5267] = 80'h00000000000000000000;
mem[5268] = 80'h00000000000000000000;
mem[5269] = 80'h00000000000000000000;
mem[5270] = 80'h10100000010000010010;
mem[5271] = 80'h00109400000208004500;
mem[5272] = 80'h0010002f60d90000fffd;
mem[5273] = 80'h0010d89fc0550102c000;
mem[5274] = 80'h00100001ffabffabffab;
mem[5275] = 80'h0010ff26275788a497f4;
mem[5276] = 80'h0010d376d3b866a515c2;
mem[5277] = 80'h00103a73d0de891bac87;
mem[5278] = 80'h01112500000000000000;
mem[5279] = 80'h00000000000000000000;
mem[5280] = 80'h10100000010000010010;
mem[5281] = 80'h00109400000208004500;
mem[5282] = 80'h0010002f60da0000fffd;
mem[5283] = 80'h0010d89ec0550102c000;
mem[5284] = 80'h00100001ffabffabffab;
mem[5285] = 80'h0010ff25b535fdcc1db3;
mem[5286] = 80'h0010132aa43050bb6489;
mem[5287] = 80'h0010c817a96d510a999e;
mem[5288] = 80'h01116800000000000000;
mem[5289] = 80'h00000000000000000000;
mem[5290] = 80'h00000000000000000000;
mem[5291] = 80'h00000000000000000000;
mem[5292] = 80'h10100000010000010010;
mem[5293] = 80'h00109400000208004500;
mem[5294] = 80'h0010002f60db0000fffd;
mem[5295] = 80'h0010d89dc0550102c000;
mem[5296] = 80'h00100001ffabffabffab;
mem[5297] = 80'h0010ff24c4ebd1146471;
mem[5298] = 80'h0010ace176b7bd4eb4c0;
mem[5299] = 80'h001099d137ef9e9ab48d;
mem[5300] = 80'h0111e500000000000000;
mem[5301] = 80'h00000000000000000000;
mem[5302] = 80'h00000000000000000000;
mem[5303] = 80'h00000000000000000000;
mem[5304] = 80'h10100000010000010010;
mem[5305] = 80'h00109400000208004500;
mem[5306] = 80'h0010002f60dc0000fffd;
mem[5307] = 80'h0010d89cc0550102c000;
mem[5308] = 80'h00100001ffabffabffab;
mem[5309] = 80'h0010ff23e02f3bc570fe;
mem[5310] = 80'h00102c5999a6d17255f8;
mem[5311] = 80'h00107c185465b58386f7;
mem[5312] = 80'h01110d00000000000000;
mem[5313] = 80'h00000000000000000000;
mem[5314] = 80'h10100000010000010010;
mem[5315] = 80'h00109400000208004500;
mem[5316] = 80'h0010002f60dd0000fffd;
mem[5317] = 80'h0010d89bc0550102c000;
mem[5318] = 80'h00100001ffabffabffab;
mem[5319] = 80'h0010ff2291f1171d093c;
mem[5320] = 80'h001093924b213c878581;
mem[5321] = 80'h00102ddb5ffb1f8ab667;
mem[5322] = 80'h0111ab00000000000000;
mem[5323] = 80'h00000000000000000000;
mem[5324] = 80'h10100000010000010010;
mem[5325] = 80'h00109400000208004500;
mem[5326] = 80'h0010002f60de0000fffd;
mem[5327] = 80'h0010d89ac0550102c000;
mem[5328] = 80'h00100001ffabffabffab;
mem[5329] = 80'h0010ff2103936275837b;
mem[5330] = 80'h001053ce3ca90a99f50a;
mem[5331] = 80'h0010df9e42a0648ab6c9;
mem[5332] = 80'h0111df00000000000000;
mem[5333] = 80'h00000000000000000000;
mem[5334] = 80'h00000000000000000000;
mem[5335] = 80'h00000000000000000000;
mem[5336] = 80'h00000000000000000000;
mem[5337] = 80'h10100000010000010010;
mem[5338] = 80'h00109400000208004500;
mem[5339] = 80'h0010002f60df0000fffd;
mem[5340] = 80'h0010d899c0550102c000;
mem[5341] = 80'h00100001ffabffabffab;
mem[5342] = 80'h0010ff20724d4eadfab9;
mem[5343] = 80'h0010ec05ee2ee76c2583;
mem[5344] = 80'h00108e4e88b7461beb78;
mem[5345] = 80'h01118f00000000000000;
mem[5346] = 80'h00000000000000000000;
mem[5347] = 80'h10100000010000010010;
mem[5348] = 80'h00109400000208004500;
mem[5349] = 80'h0010002f60e00000fffd;
mem[5350] = 80'h0010d898c0550102c000;
mem[5351] = 80'h00100001ffabffabffab;
mem[5352] = 80'h0010ff1f0170de2c3388;
mem[5353] = 80'h0010d6b1ab3207421e62;
mem[5354] = 80'h0010159194a19b76b9b9;
mem[5355] = 80'h0111e900000000000000;
mem[5356] = 80'h00000000000000000000;
mem[5357] = 80'h00000000000000000000;
mem[5358] = 80'h00000000000000000000;
mem[5359] = 80'h10100000010000010010;
mem[5360] = 80'h00109400000208004500;
mem[5361] = 80'h0010002f60e10000fffd;
mem[5362] = 80'h0010d897c0550102c000;
mem[5363] = 80'h00100001ffabffabffab;
mem[5364] = 80'h0010ff1e70aef2f44a4a;
mem[5365] = 80'h0010697a79b5eab7ce7b;
mem[5366] = 80'h00104459b536bce8376d;
mem[5367] = 80'h01119700000000000000;
mem[5368] = 80'h00000000000000000000;
mem[5369] = 80'h10100000010000010010;
mem[5370] = 80'h00109400000208004500;
mem[5371] = 80'h0010002f60e20000fffd;
mem[5372] = 80'h0010d896c0550102c000;
mem[5373] = 80'h00100001ffabffabffab;
mem[5374] = 80'h0010ff1de2cc879cc00d;
mem[5375] = 80'h0010a9260e3ddca9bef1;
mem[5376] = 80'h0010b62f993c33b566d8;
mem[5377] = 80'h0111f600000000000000;
mem[5378] = 80'h00000000000000000000;
mem[5379] = 80'h00000000000000000000;
mem[5380] = 80'h00000000000000000000;
mem[5381] = 80'h10100000010000010010;
mem[5382] = 80'h00109400000208004500;
mem[5383] = 80'h0010002f60e30000fffd;
mem[5384] = 80'h0010d895c0550102c000;
mem[5385] = 80'h00100001ffabffabffab;
mem[5386] = 80'h0010ff1c9312ab44b9cf;
mem[5387] = 80'h001016eddcba315c6978;
mem[5388] = 80'h0010e77ac3c4ce35dbd0;
mem[5389] = 80'h01118b00000000000000;
mem[5390] = 80'h00000000000000000000;
mem[5391] = 80'h10100000010000010010;
mem[5392] = 80'h00109400000208004500;
mem[5393] = 80'h0010002f60e40000fffd;
mem[5394] = 80'h0010d894c0550102c000;
mem[5395] = 80'h00100001ffabffabffab;
mem[5396] = 80'h0010ff1bb7d64195ad40;
mem[5397] = 80'h0010965533ab5d608803;
mem[5398] = 80'h001002eb3fe8670db07b;
mem[5399] = 80'h0111e900000000000000;
mem[5400] = 80'h00000000000000000000;
mem[5401] = 80'h00000000000000000000;
mem[5402] = 80'h00000000000000000000;
mem[5403] = 80'h10100000010000010010;
mem[5404] = 80'h00109400000208004500;
mem[5405] = 80'h0010002f60e50000fffd;
mem[5406] = 80'h0010d893c0550102c000;
mem[5407] = 80'h00100001ffabffabffab;
mem[5408] = 80'h0010ff1ac6086d4dd482;
mem[5409] = 80'h0010299ee12cb095587a;
mem[5410] = 80'h0010532834095d797643;
mem[5411] = 80'h01111700000000000000;
mem[5412] = 80'h00000000000000000000;
mem[5413] = 80'h10100000010000010010;
mem[5414] = 80'h00109400000208004500;
mem[5415] = 80'h0010002f60e60000fffd;
mem[5416] = 80'h0010d892c0550102c000;
mem[5417] = 80'h00100001ffabffabffab;
mem[5418] = 80'h0010ff19546a18255ec5;
mem[5419] = 80'h0010e9c296a4868b28b1;
mem[5420] = 80'h0010a160e58c7ebbfa61;
mem[5421] = 80'h01117c00000000000000;
mem[5422] = 80'h00000000000000000000;
mem[5423] = 80'h00000000000000000000;
mem[5424] = 80'h00000000000000000000;
mem[5425] = 80'h10100000010000010010;
mem[5426] = 80'h00109400000208004500;
mem[5427] = 80'h0010002f60e70000fffd;
mem[5428] = 80'h0010d891c0550102c000;
mem[5429] = 80'h00100001ffabffabffab;
mem[5430] = 80'h0010ff1825b434fd2707;
mem[5431] = 80'h0010560944236b7ef8f8;
mem[5432] = 80'h0010f0a67be413890e3b;
mem[5433] = 80'h01116d00000000000000;
mem[5434] = 80'h00000000000000000000;
mem[5435] = 80'h10100000010000010010;
mem[5436] = 80'h00109400000208004500;
mem[5437] = 80'h0010002f60e80000fffd;
mem[5438] = 80'h0010d890c0550102c000;
mem[5439] = 80'h00100001ffabffabffab;
mem[5440] = 80'h0010ff171de3cd8777da;
mem[5441] = 80'h0010e8b348865ef2eac1;
mem[5442] = 80'h00106ac112f3a4a808a0;
mem[5443] = 80'h01110300000000000000;
mem[5444] = 80'h00000000000000000000;
mem[5445] = 80'h10100000010000010010;
mem[5446] = 80'h00109400000208004500;
mem[5447] = 80'h0010002f60e90000fffd;
mem[5448] = 80'h0010d88fc0550102c000;
mem[5449] = 80'h00100001ffabffabffab;
mem[5450] = 80'h0010ff166c3de15f0e18;
mem[5451] = 80'h001057789a01b3073a80;
mem[5452] = 80'h00103b8e25a464259f59;
mem[5453] = 80'h0111e100000000000000;
mem[5454] = 80'h00000000000000000000;
mem[5455] = 80'h00000000000000000000;
mem[5456] = 80'h00000000000000000000;
mem[5457] = 80'h10100000010000010010;
mem[5458] = 80'h00109400000208004500;
mem[5459] = 80'h0010002f60ea0000fffd;
mem[5460] = 80'h0010d88ec0550102c000;
mem[5461] = 80'h00100001ffabffabffab;
mem[5462] = 80'h0010ff15fe5f9437845f;
mem[5463] = 80'h00109724ed8985194a53;
mem[5464] = 80'h0010c94c2e8b9d011aea;
mem[5465] = 80'h01115500000000000000;
mem[5466] = 80'h00000000000000000000;
mem[5467] = 80'h00000000000000000000;
mem[5468] = 80'h00000000000000000000;
mem[5469] = 80'h10100000010000010010;
mem[5470] = 80'h00109400000208004500;
mem[5471] = 80'h0010002f60eb0000fffd;
mem[5472] = 80'h0010d88dc0550102c000;
mem[5473] = 80'h00100001ffabffabffab;
mem[5474] = 80'h0010ff148f81b8effd9d;
mem[5475] = 80'h001028ef3f0e68ec9a12;
mem[5476] = 80'h0010980319dc9dd9c4c6;
mem[5477] = 80'h01118500000000000000;
mem[5478] = 80'h10100000010000010010;
mem[5479] = 80'h00109400000208004500;
mem[5480] = 80'h0010002f60ec0000fffd;
mem[5481] = 80'h0010d88cc0550102c000;
mem[5482] = 80'h00100001ffabffabffab;
mem[5483] = 80'h0010ff13ab45523ee912;
mem[5484] = 80'h0010a857d01f04d07aa1;
mem[5485] = 80'h00107d3a28327c1b70c2;
mem[5486] = 80'h01112c00000000000000;
mem[5487] = 80'h00000000000000000000;
mem[5488] = 80'h00000000000000000000;
mem[5489] = 80'h00000000000000000000;
mem[5490] = 80'h10100000010000010010;
mem[5491] = 80'h00109400000208004500;
mem[5492] = 80'h0010002f60ed0000fffd;
mem[5493] = 80'h0010d88bc0550102c000;
mem[5494] = 80'h00100001ffabffabffab;
mem[5495] = 80'h0010ff12da9b7ee690d0;
mem[5496] = 80'h0010179c0298e925aae0;
mem[5497] = 80'h00102c751feb1b6ab768;
mem[5498] = 80'h0111b200000000000000;
mem[5499] = 80'h00000000000000000000;
mem[5500] = 80'h10100000010000010010;
mem[5501] = 80'h00109400000208004500;
mem[5502] = 80'h0010002f60ee0000fffd;
mem[5503] = 80'h0010d88ac0550102c000;
mem[5504] = 80'h00100001ffabffabffab;
mem[5505] = 80'h0010ff1148f90b8e1a97;
mem[5506] = 80'h0010d7c07510df3bda53;
mem[5507] = 80'h0010debc3eb26de23996;
mem[5508] = 80'h0111e800000000000000;
mem[5509] = 80'h00000000000000000000;
mem[5510] = 80'h00000000000000000000;
mem[5511] = 80'h00000000000000000000;
mem[5512] = 80'h10100000010000010010;
mem[5513] = 80'h00109400000208004500;
mem[5514] = 80'h0010002f60ef0000fffd;
mem[5515] = 80'h0010d889c0550102c000;
mem[5516] = 80'h00100001ffabffabffab;
mem[5517] = 80'h0010ff10392727566355;
mem[5518] = 80'h0010680ba79732ce0a53;
mem[5519] = 80'h00108fcdf48a6bbf8350;
mem[5520] = 80'h01115a00000000000000;
mem[5521] = 80'h00000000000000000000;
mem[5522] = 80'h10100000010000010010;
mem[5523] = 80'h00109400000208004500;
mem[5524] = 80'h0010002f60f00000fffd;
mem[5525] = 80'h0010d888c0550102c000;
mem[5526] = 80'h00100001ffabffabffab;
mem[5527] = 80'h0010ff0f3856f97abb2c;
mem[5528] = 80'h0010aab46c5ab423ffaf;
mem[5529] = 80'h0010ea4e7ac0e39605aa;
mem[5530] = 80'h0111a200000000000000;
mem[5531] = 80'h00000000000000000000;
mem[5532] = 80'h00000000000000000000;
mem[5533] = 80'h00000000000000000000;
mem[5534] = 80'h00000000000000000000;
mem[5535] = 80'h10100000010000010010;
mem[5536] = 80'h00109400000208004500;
mem[5537] = 80'h0010002f60f10000fffd;
mem[5538] = 80'h0010d887c0550102c000;
mem[5539] = 80'h00100001ffabffabffab;
mem[5540] = 80'h0010ff0e4988d5a2c2ee;
mem[5541] = 80'h0010157fbedd59d62f2e;
mem[5542] = 80'h0010bb17195eecfad3de;
mem[5543] = 80'h0111bf00000000000000;
mem[5544] = 80'h10100000010000010010;
mem[5545] = 80'h00109400000208004500;
mem[5546] = 80'h0010002f60f20000fffd;
mem[5547] = 80'h0010d886c0550102c000;
mem[5548] = 80'h00100001ffabffabffab;
mem[5549] = 80'h0010ff0ddbeaa0ca48a9;
mem[5550] = 80'h0010d523c9556fc85fbd;
mem[5551] = 80'h001049d8debba4955799;
mem[5552] = 80'h0111e300000000000000;
mem[5553] = 80'h00000000000000000000;
mem[5554] = 80'h00000000000000000000;
mem[5555] = 80'h00000000000000000000;
mem[5556] = 80'h10100000010000010010;
mem[5557] = 80'h00109400000208004500;
mem[5558] = 80'h0010002f60f30000fffd;
mem[5559] = 80'h0010d885c0550102c000;
mem[5560] = 80'h00100001ffabffabffab;
mem[5561] = 80'h0010ff0caa348c12316b;
mem[5562] = 80'h00106ae81bd2823d8fbc;
mem[5563] = 80'h0010189a25f2c1d09eab;
mem[5564] = 80'h0111bf00000000000000;
mem[5565] = 80'h00000000000000000000;
mem[5566] = 80'h10100000010000010010;
mem[5567] = 80'h00109400000208004500;
mem[5568] = 80'h0010002f60f40000fffd;
mem[5569] = 80'h0010d884c0550102c000;
mem[5570] = 80'h00100001ffabffabffab;
mem[5571] = 80'h0010ff0b8ef066c325e4;
mem[5572] = 80'h0010ea50f4c3ee016ecf;
mem[5573] = 80'h0010fd8270f33aec82e4;
mem[5574] = 80'h0111d200000000000000;
mem[5575] = 80'h00000000000000000000;
mem[5576] = 80'h00000000000000000000;
mem[5577] = 80'h00000000000000000000;
mem[5578] = 80'h10100000010000010010;
mem[5579] = 80'h00109400000208004500;
mem[5580] = 80'h0010002f60f50000fffd;
mem[5581] = 80'h0010d883c0550102c000;
mem[5582] = 80'h00100001ffabffabffab;
mem[5583] = 80'h0010ff0aff2e4a1b5c26;
mem[5584] = 80'h0010559b264403f4bd4d;
mem[5585] = 80'h0010acd7108c60aaebb8;
mem[5586] = 80'h01111c00000000000000;
mem[5587] = 80'h00000000000000000000;
mem[5588] = 80'h10100000010000010010;
mem[5589] = 80'h00109400000208004500;
mem[5590] = 80'h0010002f60f60000fffd;
mem[5591] = 80'h0010d882c0550102c000;
mem[5592] = 80'h00100001ffabffabffab;
mem[5593] = 80'h0010ff096d4c3f73d661;
mem[5594] = 80'h001095c751cc35eacdfe;
mem[5595] = 80'h00105e1e313a027c5e7a;
mem[5596] = 80'h01118500000000000000;
mem[5597] = 80'h00000000000000000000;
mem[5598] = 80'h00000000000000000000;
mem[5599] = 80'h00000000000000000000;
mem[5600] = 80'h00000000000000000000;
mem[5601] = 80'h10100000010000010010;
mem[5602] = 80'h00109400000208004500;
mem[5603] = 80'h0010002f60f70000fffd;
mem[5604] = 80'h0010d881c0550102c000;
mem[5605] = 80'h00100001ffabffabffab;
mem[5606] = 80'h0010ff081c9213abafa3;
mem[5607] = 80'h00102a0c834bd81f1dbf;
mem[5608] = 80'h00100f51068f671d84c6;
mem[5609] = 80'h01110400000000000000;
mem[5610] = 80'h10100000010000010010;
mem[5611] = 80'h00109400000208004500;
mem[5612] = 80'h0010002f60f80000fffd;
mem[5613] = 80'h0010d880c0550102c000;
mem[5614] = 80'h00100001ffabffabffab;
mem[5615] = 80'h0010ff0724c5ead1ff7e;
mem[5616] = 80'h001094b68feeed930f09;
mem[5617] = 80'h0010953dc96271ab18cd;
mem[5618] = 80'h0111c000000000000000;
mem[5619] = 80'h00000000000000000000;
mem[5620] = 80'h00000000000000000000;
mem[5621] = 80'h00000000000000000000;
mem[5622] = 80'h10100000010000010010;
mem[5623] = 80'h00109400000208004500;
mem[5624] = 80'h0010002f60f90000fffd;
mem[5625] = 80'h0010d87fc0550102c000;
mem[5626] = 80'h00100001ffabffabffab;
mem[5627] = 80'h0010ff06551bc60986bc;
mem[5628] = 80'h00102b7d5d690066df48;
mem[5629] = 80'h0010c472fe0f33bcfff0;
mem[5630] = 80'h01114900000000000000;
mem[5631] = 80'h00000000000000000000;
mem[5632] = 80'h10100000010000010010;
mem[5633] = 80'h00109400000208004500;
mem[5634] = 80'h0010002f60fa0000fffd;
mem[5635] = 80'h0010d87ec0550102c000;
mem[5636] = 80'h00100001ffabffabffab;
mem[5637] = 80'h0010ff05c779b3610cfb;
mem[5638] = 80'h0010eb212ae13678af1b;
mem[5639] = 80'h001036ab6de1d8d1c0b3;
mem[5640] = 80'h0111b600000000000000;
mem[5641] = 80'h00000000000000000000;
mem[5642] = 80'h00000000000000000000;
mem[5643] = 80'h00000000000000000000;
mem[5644] = 80'h10100000010000010010;
mem[5645] = 80'h00109400000208004500;
mem[5646] = 80'h0010002f60fb0000fffd;
mem[5647] = 80'h0010d87dc0550102c000;
mem[5648] = 80'h00100001ffabffabffab;
mem[5649] = 80'h0010ff04b6a79fb97539;
mem[5650] = 80'h001054eaf866db8d7f5b;
mem[5651] = 80'h001067d76b4eb93f2f24;
mem[5652] = 80'h01118c00000000000000;
mem[5653] = 80'h00000000000000000000;
mem[5654] = 80'h00000000000000000000;
mem[5655] = 80'h00000000000000000000;
mem[5656] = 80'h10100000010000010010;
mem[5657] = 80'h00109400000208004500;
mem[5658] = 80'h0010002f60fc0000fffd;
mem[5659] = 80'h0010d87cc0550102c000;
mem[5660] = 80'h00100001ffabffabffab;
mem[5661] = 80'h0010ff039263756861b6;
mem[5662] = 80'h0010d4521777b7b19e68;
mem[5663] = 80'h001082c2f2d2df3895bd;
mem[5664] = 80'h0111ce00000000000000;
mem[5665] = 80'h00000000000000000000;
mem[5666] = 80'h10100000010000010010;
mem[5667] = 80'h00109400000208004500;
mem[5668] = 80'h0010002f60fd0000fffd;
mem[5669] = 80'h0010d87bc0550102c000;
mem[5670] = 80'h00100001ffabffabffab;
mem[5671] = 80'h0010ff02e3bd59b01874;
mem[5672] = 80'h00106b99c5f05a444e29;
mem[5673] = 80'h0010d38dc595376c6bd2;
mem[5674] = 80'h0111c200000000000000;
mem[5675] = 80'h00000000000000000000;
mem[5676] = 80'h10100000010000010010;
mem[5677] = 80'h00109400000208004500;
mem[5678] = 80'h0010002f60fe0000fffd;
mem[5679] = 80'h0010d87ac0550102c000;
mem[5680] = 80'h00100001ffabffabffab;
mem[5681] = 80'h0010ff0171df2cd89233;
mem[5682] = 80'h0010abc5b2786c5a3e9a;
mem[5683] = 80'h00102144e49bc0c19d69;
mem[5684] = 80'h0111f700000000000000;
mem[5685] = 80'h00000000000000000000;
mem[5686] = 80'h00000000000000000000;
mem[5687] = 80'h00000000000000000000;
mem[5688] = 80'h00000000000000000000;
mem[5689] = 80'h10100000010000010010;
mem[5690] = 80'h00109400000208004500;
mem[5691] = 80'h0010002f60ff0000fffd;
mem[5692] = 80'h0010d879c0550102c000;
mem[5693] = 80'h00100001ffabffabffab;
mem[5694] = 80'h0010ff0000010000ebf1;
mem[5695] = 80'h0010140e60ff81afef1b;
mem[5696] = 80'h0010702ab70907a68907;
mem[5697] = 80'h01117400000000000000;
mem[5698] = 80'h00000000000000000000;
mem[5699] = 80'h10100000010000010010;
mem[5700] = 80'h00109400000208004500;
mem[5701] = 80'h0010002f61000000fffd;
mem[5702] = 80'h0010d878c0550102c000;
mem[5703] = 80'h00100001ffabffabffab;
mem[5704] = 80'h0010ffff2f4b1bb73cb0;
mem[5705] = 80'h00108148d082dafca0eb;
mem[5706] = 80'h0010bfca2fcfbafdbb45;
mem[5707] = 80'h01119e00000000000000;
mem[5708] = 80'h00000000000000000000;
mem[5709] = 80'h00000000000000000000;
mem[5710] = 80'h00000000000000000000;
mem[5711] = 80'h10100000010000010010;
mem[5712] = 80'h00109400000208004500;
mem[5713] = 80'h0010002f61010000fffd;
mem[5714] = 80'h0010d877c0550102c000;
mem[5715] = 80'h00100001ffabffabffab;
mem[5716] = 80'h0010fffe5e95376f4572;
mem[5717] = 80'h00103e830205370970ed;
mem[5718] = 80'h0010ee1143fa09f9eaac;
mem[5719] = 80'h01114300000000000000;
mem[5720] = 80'h00000000000000000000;
mem[5721] = 80'h10100000010000010010;
mem[5722] = 80'h00109400000208004500;
mem[5723] = 80'h0010002f61020000fffd;
mem[5724] = 80'h0010d876c0550102c000;
mem[5725] = 80'h00100001ffabffabffab;
mem[5726] = 80'h0010fffdccf74207cf35;
mem[5727] = 80'h0010fedf758d01170066;
mem[5728] = 80'h00101c545e8f3069c3d7;
mem[5729] = 80'h0111a400000000000000;
mem[5730] = 80'h00000000000000000000;
mem[5731] = 80'h00000000000000000000;
mem[5732] = 80'h00000000000000000000;
mem[5733] = 80'h10100000010000010010;
mem[5734] = 80'h00109400000208004500;
mem[5735] = 80'h0010002f61030000fffd;
mem[5736] = 80'h0010d875c0550102c000;
mem[5737] = 80'h00100001ffabffabffab;
mem[5738] = 80'h0010fffcbd296edfb6f7;
mem[5739] = 80'h00104114a70aece2d0ff;
mem[5740] = 80'h00104d87e779416727b5;
mem[5741] = 80'h01110600000000000000;
mem[5742] = 80'h00000000000000000000;
mem[5743] = 80'h10100000010000010010;
mem[5744] = 80'h00109400000208004500;
mem[5745] = 80'h0010002f61040000fffd;
mem[5746] = 80'h0010d874c0550102c000;
mem[5747] = 80'h00100001ffabffabffab;
mem[5748] = 80'h0010fffb99ed840ea278;
mem[5749] = 80'h0010c1ac481b80de3184;
mem[5750] = 80'h0010a8161b4ebf924327;
mem[5751] = 80'h01113800000000000000;
mem[5752] = 80'h00000000000000000000;
mem[5753] = 80'h00000000000000000000;
mem[5754] = 80'h00000000000000000000;
mem[5755] = 80'h10100000010000010010;
mem[5756] = 80'h00109400000208004500;
mem[5757] = 80'h0010002f61050000fffd;
mem[5758] = 80'h0010d873c0550102c000;
mem[5759] = 80'h00100001ffabffabffab;
mem[5760] = 80'h0010fffae833a8d6dbba;
mem[5761] = 80'h00107e679a9c6d2be18d;
mem[5762] = 80'h0010f9dd49a4e7486cac;
mem[5763] = 80'h01112b00000000000000;
mem[5764] = 80'h00000000000000000000;
mem[5765] = 80'h10100000010000010010;
mem[5766] = 80'h00109400000208004500;
mem[5767] = 80'h0010002f61060000fffd;
mem[5768] = 80'h0010d872c0550102c000;
mem[5769] = 80'h00100001ffabffabffab;
mem[5770] = 80'h0010fff97a51ddbe51fd;
mem[5771] = 80'h0010be3bed145b359106;
mem[5772] = 80'h00100b9854d45d076311;
mem[5773] = 80'h0111c500000000000000;
mem[5774] = 80'h00000000000000000000;
mem[5775] = 80'h00000000000000000000;
mem[5776] = 80'h00000000000000000000;
mem[5777] = 80'h10100000010000010010;
mem[5778] = 80'h00109400000208004500;
mem[5779] = 80'h0010002f61070000fffd;
mem[5780] = 80'h0010d871c0550102c000;
mem[5781] = 80'h00100001ffabffabffab;
mem[5782] = 80'h0010fff80b8ff166283f;
mem[5783] = 80'h001001f03f93b6c0417f;
mem[5784] = 80'h00105a5b5fb3e69f711f;
mem[5785] = 80'h0111f400000000000000;
mem[5786] = 80'h00000000000000000000;
mem[5787] = 80'h10100000010000010010;
mem[5788] = 80'h00109400000208004500;
mem[5789] = 80'h0010002f61080000fffd;
mem[5790] = 80'h0010d870c0550102c000;
mem[5791] = 80'h00100001ffabffabffab;
mem[5792] = 80'h0010fff733d8081c78e2;
mem[5793] = 80'h0010bf4a3336834c4c40;
mem[5794] = 80'h0010c0f9c22a05949d13;
mem[5795] = 80'h0111e700000000000000;
mem[5796] = 80'h00000000000000000000;
mem[5797] = 80'h10100000010000010010;
mem[5798] = 80'h00109400000208004500;
mem[5799] = 80'h0010002f61090000fffd;
mem[5800] = 80'h0010d86fc0550102c000;
mem[5801] = 80'h00100001ffabffabffab;
mem[5802] = 80'h0010fff6420624c40120;
mem[5803] = 80'h00100081e1b16eb99c09;
mem[5804] = 80'h0010913f5ce9bcac91b5;
mem[5805] = 80'h01119300000000000000;
mem[5806] = 80'h00000000000000000000;
mem[5807] = 80'h00000000000000000000;
mem[5808] = 80'h00000000000000000000;
mem[5809] = 80'h10100000010000010010;
mem[5810] = 80'h00109400000208004500;
mem[5811] = 80'h0010002f610a0000fffd;
mem[5812] = 80'h0010d86ec0550102c000;
mem[5813] = 80'h00100001ffabffabffab;
mem[5814] = 80'h0010fff5d06451ac8b67;
mem[5815] = 80'h0010c0dd963958a7ecc2;
mem[5816] = 80'h001063778d98c4abb1fe;
mem[5817] = 80'h01117400000000000000;
mem[5818] = 80'h00000000000000000000;
mem[5819] = 80'h00000000000000000000;
mem[5820] = 80'h00000000000000000000;
mem[5821] = 80'h10100000010000010010;
mem[5822] = 80'h00109400000208004500;
mem[5823] = 80'h0010002f610b0000fffd;
mem[5824] = 80'h0010d86dc0550102c000;
mem[5825] = 80'h00100001ffabffabffab;
mem[5826] = 80'h0010fff4a1ba7d74f2a5;
mem[5827] = 80'h00107f1644beb5523c9b;
mem[5828] = 80'h001032b260c1a4ea459c;
mem[5829] = 80'h01119a00000000000000;
mem[5830] = 80'h10100000010000010010;
mem[5831] = 80'h00109400000208004500;
mem[5832] = 80'h0010002f610c0000fffd;
mem[5833] = 80'h0010d86cc0550102c000;
mem[5834] = 80'h00100001ffabffabffab;
mem[5835] = 80'h0010fff3857e97a5e62a;
mem[5836] = 80'h0010ffaeabafd96edd20;
mem[5837] = 80'h0010d735c898fa455489;
mem[5838] = 80'h01118600000000000000;
mem[5839] = 80'h00000000000000000000;
mem[5840] = 80'h00000000000000000000;
mem[5841] = 80'h00000000000000000000;
mem[5842] = 80'h10100000010000010010;
mem[5843] = 80'h00109400000208004500;
mem[5844] = 80'h0010002f610d0000fffd;
mem[5845] = 80'h0010d86bc0550102c000;
mem[5846] = 80'h00100001ffabffabffab;
mem[5847] = 80'h0010fff2f4a0bb7d9fe8;
mem[5848] = 80'h001040657928349b0d69;
mem[5849] = 80'h001086f35680d610f067;
mem[5850] = 80'h01118100000000000000;
mem[5851] = 80'h00000000000000000000;
mem[5852] = 80'h10100000010000010010;
mem[5853] = 80'h00109400000208004500;
mem[5854] = 80'h0010002f610e0000fffd;
mem[5855] = 80'h0010d86ac0550102c000;
mem[5856] = 80'h00100001ffabffabffab;
mem[5857] = 80'h0010fff166c2ce1515af;
mem[5858] = 80'h001080390ea002857da1;
mem[5859] = 80'h001074eed4985c1e8e1d;
mem[5860] = 80'h01119500000000000000;
mem[5861] = 80'h00000000000000000000;
mem[5862] = 80'h00000000000000000000;
mem[5863] = 80'h00000000000000000000;
mem[5864] = 80'h10100000010000010010;
mem[5865] = 80'h00109400000208004500;
mem[5866] = 80'h0010002f610f0000fffd;
mem[5867] = 80'h0010d869c0550102c000;
mem[5868] = 80'h00100001ffabffabffab;
mem[5869] = 80'h0010fff0171ce2cd6c6d;
mem[5870] = 80'h00103ff2dc27ef70add8;
mem[5871] = 80'h0010252ddf26db579e86;
mem[5872] = 80'h0111db00000000000000;
mem[5873] = 80'h00000000000000000000;
mem[5874] = 80'h10100000010000010010;
mem[5875] = 80'h00109400000208004500;
mem[5876] = 80'h0010002f61100000fffd;
mem[5877] = 80'h0010d868c0550102c000;
mem[5878] = 80'h00100001ffabffabffab;
mem[5879] = 80'h0010ffef166d3ce1b414;
mem[5880] = 80'h0010fd4d17ea699d582c;
mem[5881] = 80'h00104027f883e86a8082;
mem[5882] = 80'h01110c00000000000000;
mem[5883] = 80'h00000000000000000000;
mem[5884] = 80'h00000000000000000000;
mem[5885] = 80'h00000000000000000000;
mem[5886] = 80'h00000000000000000000;
mem[5887] = 80'h10100000010000010010;
mem[5888] = 80'h00109400000208004500;
mem[5889] = 80'h0010002f61110000fffd;
mem[5890] = 80'h0010d867c0550102c000;
mem[5891] = 80'h00100001ffabffabffab;
mem[5892] = 80'h0010ffee67b31039cdd6;
mem[5893] = 80'h00104286c56d846889a5;
mem[5894] = 80'h001011c0028c8f38378e;
mem[5895] = 80'h01117f00000000000000;
mem[5896] = 80'h10100000010000010010;
mem[5897] = 80'h00109400000208004500;
mem[5898] = 80'h0010002f61120000fffd;
mem[5899] = 80'h0010d866c0550102c000;
mem[5900] = 80'h00100001ffabffabffab;
mem[5901] = 80'h0010ffedf5d165514791;
mem[5902] = 80'h001082dab2e5b276f92e;
mem[5903] = 80'h0010e3851f72789fb05e;
mem[5904] = 80'h01113c00000000000000;
mem[5905] = 80'h00000000000000000000;
mem[5906] = 80'h00000000000000000000;
mem[5907] = 80'h00000000000000000000;
mem[5908] = 80'h10100000010000010010;
mem[5909] = 80'h00109400000208004500;
mem[5910] = 80'h0010002f61130000fffd;
mem[5911] = 80'h0010d865c0550102c000;
mem[5912] = 80'h00100001ffabffabffab;
mem[5913] = 80'h0010ffec840f49893e53;
mem[5914] = 80'h00103d1160625f832937;
mem[5915] = 80'h0010b24d3eabdca96731;
mem[5916] = 80'h01111000000000000000;
mem[5917] = 80'h00000000000000000000;
mem[5918] = 80'h10100000010000010010;
mem[5919] = 80'h00109400000208004500;
mem[5920] = 80'h0010002f61140000fffd;
mem[5921] = 80'h0010d864c0550102c000;
mem[5922] = 80'h00100001ffabffabffab;
mem[5923] = 80'h0010ffeba0cba3582adc;
mem[5924] = 80'h0010bda98f7333bfc84d;
mem[5925] = 80'h001057eff3f9fb83fd4d;
mem[5926] = 80'h0111c500000000000000;
mem[5927] = 80'h00000000000000000000;
mem[5928] = 80'h00000000000000000000;
mem[5929] = 80'h00000000000000000000;
mem[5930] = 80'h10100000010000010010;
mem[5931] = 80'h00109400000208004500;
mem[5932] = 80'h0010002f61150000fffd;
mem[5933] = 80'h0010d863c0550102c000;
mem[5934] = 80'h00100001ffabffabffab;
mem[5935] = 80'h0010ffead1158f80531e;
mem[5936] = 80'h001002625df4de4a18c4;
mem[5937] = 80'h0010063f39bcb4b6da22;
mem[5938] = 80'h01111600000000000000;
mem[5939] = 80'h00000000000000000000;
mem[5940] = 80'h10100000010000010010;
mem[5941] = 80'h00109400000208004500;
mem[5942] = 80'h0010002f61160000fffd;
mem[5943] = 80'h0010d862c0550102c000;
mem[5944] = 80'h00100001ffabffabffab;
mem[5945] = 80'h0010ffe94377fae8d959;
mem[5946] = 80'h0010c23e2a7ce854684f;
mem[5947] = 80'h0010f47a248291a739d5;
mem[5948] = 80'h0111f600000000000000;
mem[5949] = 80'h00000000000000000000;
mem[5950] = 80'h00000000000000000000;
mem[5951] = 80'h00000000000000000000;
mem[5952] = 80'h00000000000000000000;
mem[5953] = 80'h10100000010000010010;
mem[5954] = 80'h00109400000208004500;
mem[5955] = 80'h0010002f61170000fffd;
mem[5956] = 80'h0010d861c0550102c000;
mem[5957] = 80'h00100001ffabffabffab;
mem[5958] = 80'h0010ffe832a9d630a09b;
mem[5959] = 80'h00107df5f8fb05a1b836;
mem[5960] = 80'h0010a5b92f1f4c65e659;
mem[5961] = 80'h01118d00000000000000;
mem[5962] = 80'h10100000010000010010;
mem[5963] = 80'h00109400000208004500;
mem[5964] = 80'h0010002f61180000fffd;
mem[5965] = 80'h0010d860c0550102c000;
mem[5966] = 80'h00100001ffabffabffab;
mem[5967] = 80'h0010ffe70afe2f4af046;
mem[5968] = 80'h0010c34ff45e302daa88;
mem[5969] = 80'h00103f5c49c8b95b0a53;
mem[5970] = 80'h0111ff00000000000000;
mem[5971] = 80'h00000000000000000000;
mem[5972] = 80'h00000000000000000000;
mem[5973] = 80'h00000000000000000000;
mem[5974] = 80'h10100000010000010010;
mem[5975] = 80'h00109400000208004500;
mem[5976] = 80'h0010002f61190000fffd;
mem[5977] = 80'h0010d85fc0550102c000;
mem[5978] = 80'h00100001ffabffabffab;
mem[5979] = 80'h0010ffe67b2003928984;
mem[5980] = 80'h00107c8426d9ddd87ac1;
mem[5981] = 80'h00106e9ad74fb5980918;
mem[5982] = 80'h0111bd00000000000000;
mem[5983] = 80'h00000000000000000000;
mem[5984] = 80'h10100000010000010010;
mem[5985] = 80'h00109400000208004500;
mem[5986] = 80'h0010002f611a0000fffd;
mem[5987] = 80'h0010d85ec0550102c000;
mem[5988] = 80'h00100001ffabffabffab;
mem[5989] = 80'h0010ffe5e94276fa03c3;
mem[5990] = 80'h0010bcd85151ebc6098d;
mem[5991] = 80'h00109c095992a25bcf04;
mem[5992] = 80'h01112100000000000000;
mem[5993] = 80'h00000000000000000000;
mem[5994] = 80'h00000000000000000000;
mem[5995] = 80'h00000000000000000000;
mem[5996] = 80'h10100000010000010010;
mem[5997] = 80'h00109400000208004500;
mem[5998] = 80'h0010002f611b0000fffd;
mem[5999] = 80'h0010d85dc0550102c000;
mem[6000] = 80'h00100001ffabffabffab;
mem[6001] = 80'h0010ffe4989c5a227a01;
mem[6002] = 80'h0010031383d60633d9cc;
mem[6003] = 80'h0010cd466e2af078ceab;
mem[6004] = 80'h0111ad00000000000000;
mem[6005] = 80'h00000000000000000000;
mem[6006] = 80'h00000000000000000000;
mem[6007] = 80'h00000000000000000000;
mem[6008] = 80'h10100000010000010010;
mem[6009] = 80'h00109400000208004500;
mem[6010] = 80'h0010002f611c0000fffd;
mem[6011] = 80'h0010d85cc0550102c000;
mem[6012] = 80'h00100001ffabffabffab;
mem[6013] = 80'h0010ffe3bc58b0f36e8e;
mem[6014] = 80'h001083ab6cc76a0f38ef;
mem[6015] = 80'h00102850847fe3b7e6b1;
mem[6016] = 80'h01119200000000000000;
mem[6017] = 80'h00000000000000000000;
mem[6018] = 80'h10100000010000010010;
mem[6019] = 80'h00109400000208004500;
mem[6020] = 80'h0010002f611d0000fffd;
mem[6021] = 80'h0010d85bc0550102c000;
mem[6022] = 80'h00100001ffabffabffab;
mem[6023] = 80'h0010ffe2cd869c2b174c;
mem[6024] = 80'h00103c60be4087fae8ae;
mem[6025] = 80'h0010791fb3b4e6615153;
mem[6026] = 80'h0111d700000000000000;
mem[6027] = 80'h00000000000000000000;
mem[6028] = 80'h10100000010000010010;
mem[6029] = 80'h00109400000208004500;
mem[6030] = 80'h0010002f611e0000fffd;
mem[6031] = 80'h0010d85ac0550102c000;
mem[6032] = 80'h00100001ffabffabffab;
mem[6033] = 80'h0010ffe15fe4e9439d0b;
mem[6034] = 80'h0010fc3cc9c8b1e498ed;
mem[6035] = 80'h00108bc5534d29377544;
mem[6036] = 80'h01115600000000000000;
mem[6037] = 80'h00000000000000000000;
mem[6038] = 80'h00000000000000000000;
mem[6039] = 80'h00000000000000000000;
mem[6040] = 80'h00000000000000000000;
mem[6041] = 80'h10100000010000010010;
mem[6042] = 80'h00109400000208004500;
mem[6043] = 80'h0010002f611f0000fffd;
mem[6044] = 80'h0010d859c0550102c000;
mem[6045] = 80'h00100001ffabffabffab;
mem[6046] = 80'h0010ffe02e3ac59be4c9;
mem[6047] = 80'h001043f71b4f5c1148ac;
mem[6048] = 80'h0010da8a64f0e3279b48;
mem[6049] = 80'h01115900000000000000;
mem[6050] = 80'h00000000000000000000;
mem[6051] = 80'h10100000010000010010;
mem[6052] = 80'h00109400000208004500;
mem[6053] = 80'h0010002f61200000fffd;
mem[6054] = 80'h0010d858c0550102c000;
mem[6055] = 80'h00100001ffabffabffab;
mem[6056] = 80'h0010ffdf5d07551a2df8;
mem[6057] = 80'h001079435e53bc3f7375;
mem[6058] = 80'h001041d944e191437176;
mem[6059] = 80'h01115400000000000000;
mem[6060] = 80'h00000000000000000000;
mem[6061] = 80'h00000000000000000000;
mem[6062] = 80'h00000000000000000000;
mem[6063] = 80'h10100000010000010010;
mem[6064] = 80'h00109400000208004500;
mem[6065] = 80'h0010002f61210000fffd;
mem[6066] = 80'h0010d857c0550102c000;
mem[6067] = 80'h00100001ffabffabffab;
mem[6068] = 80'h0010ffde2cd979c2543a;
mem[6069] = 80'h0010c6888cd451caa375;
mem[6070] = 80'h001010a88e061d49918d;
mem[6071] = 80'h0111a500000000000000;
mem[6072] = 80'h00000000000000000000;
mem[6073] = 80'h10100000010000010010;
mem[6074] = 80'h00109400000208004500;
mem[6075] = 80'h0010002f61220000fffd;
mem[6076] = 80'h0010d856c0550102c000;
mem[6077] = 80'h00100001ffabffabffab;
mem[6078] = 80'h0010ffddbebb0caade7d;
mem[6079] = 80'h001006d4fb5c67d4d3f6;
mem[6080] = 80'h0010e2643addfa5ecbb2;
mem[6081] = 80'h0111b900000000000000;
mem[6082] = 80'h00000000000000000000;
mem[6083] = 80'h00000000000000000000;
mem[6084] = 80'h00000000000000000000;
mem[6085] = 80'h10100000010000010010;
mem[6086] = 80'h00109400000208004500;
mem[6087] = 80'h0010002f61230000fffd;
mem[6088] = 80'h0010d855c0550102c000;
mem[6089] = 80'h00100001ffabffabffab;
mem[6090] = 80'h0010ffdccf652072a7bf;
mem[6091] = 80'h0010b91f29db8a210277;
mem[6092] = 80'h0010b30a69eddb1f4684;
mem[6093] = 80'h0111ef00000000000000;
mem[6094] = 80'h00000000000000000000;
mem[6095] = 80'h10100000010000010010;
mem[6096] = 80'h00109400000208004500;
mem[6097] = 80'h0010002f61240000fffd;
mem[6098] = 80'h0010d854c0550102c000;
mem[6099] = 80'h00100001ffabffabffab;
mem[6100] = 80'h0010ffdbeba1caa3b330;
mem[6101] = 80'h001039a7c6cae61de314;
mem[6102] = 80'h001056114ff8263f53d2;
mem[6103] = 80'h01110200000000000000;
mem[6104] = 80'h00000000000000000000;
mem[6105] = 80'h00000000000000000000;
mem[6106] = 80'h00000000000000000000;
mem[6107] = 80'h10100000010000010010;
mem[6108] = 80'h00109400000208004500;
mem[6109] = 80'h0010002f61250000fffd;
mem[6110] = 80'h0010d853c0550102c000;
mem[6111] = 80'h00100001ffabffabffab;
mem[6112] = 80'h0010ffda9a7fe67bcaf2;
mem[6113] = 80'h0010866c144d0be83315;
mem[6114] = 80'h00100753b42d1eb22a9e;
mem[6115] = 80'h0111ae00000000000000;
mem[6116] = 80'h00000000000000000000;
mem[6117] = 80'h10100000010000010010;
mem[6118] = 80'h00109400000208004500;
mem[6119] = 80'h0010002f61260000fffd;
mem[6120] = 80'h0010d852c0550102c000;
mem[6121] = 80'h00100001ffabffabffab;
mem[6122] = 80'h0010ffd9081d931340b5;
mem[6123] = 80'h0010463063c53df64396;
mem[6124] = 80'h0010f59f001f02941372;
mem[6125] = 80'h01111700000000000000;
mem[6126] = 80'h00000000000000000000;
mem[6127] = 80'h00000000000000000000;
mem[6128] = 80'h00000000000000000000;
mem[6129] = 80'h10100000010000010010;
mem[6130] = 80'h00109400000208004500;
mem[6131] = 80'h0010002f61270000fffd;
mem[6132] = 80'h0010d851c0550102c000;
mem[6133] = 80'h00100001ffabffabffab;
mem[6134] = 80'h0010ffd879c3bfcb3977;
mem[6135] = 80'h0010f9fbb142d0039314;
mem[6136] = 80'h0010a4933036a9186e74;
mem[6137] = 80'h01112c00000000000000;
mem[6138] = 80'h00000000000000000000;
mem[6139] = 80'h10100000010000010010;
mem[6140] = 80'h00109400000208004500;
mem[6141] = 80'h0010002f61280000fffd;
mem[6142] = 80'h0010d850c0550102c000;
mem[6143] = 80'h00100001ffabffabffab;
mem[6144] = 80'h0010ffd7419446b169aa;
mem[6145] = 80'h00104741bde7e58f81d2;
mem[6146] = 80'h00103ef7a6b5bb8f4097;
mem[6147] = 80'h0111b900000000000000;
mem[6148] = 80'h00000000000000000000;
mem[6149] = 80'h10100000010000010010;
mem[6150] = 80'h00109400000208004500;
mem[6151] = 80'h0010002f61290000fffd;
mem[6152] = 80'h0010d84fc0550102c000;
mem[6153] = 80'h00100001ffabffabffab;
mem[6154] = 80'h0010ffd6304a6a691068;
mem[6155] = 80'h0010f88a6f60087a5193;
mem[6156] = 80'h00106fb8915c91525ff7;
mem[6157] = 80'h01116100000000000000;
mem[6158] = 80'h00000000000000000000;
mem[6159] = 80'h00000000000000000000;
mem[6160] = 80'h00000000000000000000;
mem[6161] = 80'h10100000010000010010;
mem[6162] = 80'h00109400000208004500;
mem[6163] = 80'h0010002f612a0000fffd;
mem[6164] = 80'h0010d84ec0550102c000;
mem[6165] = 80'h00100001ffabffabffab;
mem[6166] = 80'h0010ffd5a2281f019a2f;
mem[6167] = 80'h001038d618e83e642150;
mem[6168] = 80'h00109d79e9e46b6dec99;
mem[6169] = 80'h01113500000000000000;
mem[6170] = 80'h00000000000000000000;
mem[6171] = 80'h00000000000000000000;
mem[6172] = 80'h00000000000000000000;
mem[6173] = 80'h10100000010000010010;
mem[6174] = 80'h00109400000208004500;
mem[6175] = 80'h0010002f612b0000fffd;
mem[6176] = 80'h0010d84dc0550102c000;
mem[6177] = 80'h00100001ffabffabffab;
mem[6178] = 80'h0010ffd4d3f633d9e3ed;
mem[6179] = 80'h0010871dca6fd391f111;
mem[6180] = 80'h0010cc36de0553158328;
mem[6181] = 80'h01117f00000000000000;
mem[6182] = 80'h10100000010000010010;
mem[6183] = 80'h00109400000208004500;
mem[6184] = 80'h0010002f612c0000fffd;
mem[6185] = 80'h0010d84cc0550102c000;
mem[6186] = 80'h00100001ffabffabffab;
mem[6187] = 80'h0010ffd3f732d908f762;
mem[6188] = 80'h001007a5257ebfad17b2;
mem[6189] = 80'h001029be3c4ccd63e4d7;
mem[6190] = 80'h0111bd00000000000000;
mem[6191] = 80'h00000000000000000000;
mem[6192] = 80'h00000000000000000000;
mem[6193] = 80'h00000000000000000000;
mem[6194] = 80'h10100000010000010010;
mem[6195] = 80'h00109400000208004500;
mem[6196] = 80'h0010002f612d0000fffd;
mem[6197] = 80'h0010d84bc0550102c000;
mem[6198] = 80'h00100001ffabffabffab;
mem[6199] = 80'h0010ffd286ecf5d08ea0;
mem[6200] = 80'h0010b86ef7f95258c7f2;
mem[6201] = 80'h001078c23a5976e22e3c;
mem[6202] = 80'h0111c700000000000000;
mem[6203] = 80'h00000000000000000000;
mem[6204] = 80'h10100000010000010010;
mem[6205] = 80'h00109400000208004500;
mem[6206] = 80'h0010002f612e0000fffd;
mem[6207] = 80'h0010d84ac0550102c000;
mem[6208] = 80'h00100001ffabffabffab;
mem[6209] = 80'h0010ffd1148e80b804e7;
mem[6210] = 80'h0010783280716446b731;
mem[6211] = 80'h00108a0342e184ef1589;
mem[6212] = 80'h01119d00000000000000;
mem[6213] = 80'h00000000000000000000;
mem[6214] = 80'h00000000000000000000;
mem[6215] = 80'h00000000000000000000;
mem[6216] = 80'h10100000010000010010;
mem[6217] = 80'h00109400000208004500;
mem[6218] = 80'h0010002f612f0000fffd;
mem[6219] = 80'h0010d849c0550102c000;
mem[6220] = 80'h00100001ffabffabffab;
mem[6221] = 80'h0010ffd06550ac607d25;
mem[6222] = 80'h0010c7f952f689b36770;
mem[6223] = 80'h0010db4c75f8135baf34;
mem[6224] = 80'h01114d00000000000000;
mem[6225] = 80'h00000000000000000000;
mem[6226] = 80'h10100000010000010010;
mem[6227] = 80'h00109400000208004500;
mem[6228] = 80'h0010002f61300000fffd;
mem[6229] = 80'h0010d848c0550102c000;
mem[6230] = 80'h00100001ffabffabffab;
mem[6231] = 80'h0010ffcf6421724ca55c;
mem[6232] = 80'h00100546993b0f5e92bc;
mem[6233] = 80'h0010beca6eff15993b65;
mem[6234] = 80'h01113200000000000000;
mem[6235] = 80'h00000000000000000000;
mem[6236] = 80'h00000000000000000000;
mem[6237] = 80'h00000000000000000000;
mem[6238] = 80'h00000000000000000000;
mem[6239] = 80'h10100000010000010010;
mem[6240] = 80'h00109400000208004500;
mem[6241] = 80'h0010002f61310000fffd;
mem[6242] = 80'h0010d847c0550102c000;
mem[6243] = 80'h00100001ffabffabffab;
mem[6244] = 80'h0010ffce15ff5e94dc9e;
mem[6245] = 80'h0010ba8d4bbce2ab423d;
mem[6246] = 80'h0010ef930d388687d4d1;
mem[6247] = 80'h0111bd00000000000000;
mem[6248] = 80'h10100000010000010010;
mem[6249] = 80'h00109400000208004500;
mem[6250] = 80'h0010002f61320000fffd;
mem[6251] = 80'h0010d846c0550102c000;
mem[6252] = 80'h00100001ffabffabffab;
mem[6253] = 80'h0010ffcd879d2bfc56d9;
mem[6254] = 80'h00107ad13c34d4b532be;
mem[6255] = 80'h00101d5fb9e65f7e67f8;
mem[6256] = 80'h01111d00000000000000;
mem[6257] = 80'h00000000000000000000;
mem[6258] = 80'h00000000000000000000;
mem[6259] = 80'h00000000000000000000;
mem[6260] = 80'h10100000010000010010;
mem[6261] = 80'h00109400000208004500;
mem[6262] = 80'h0010002f61330000fffd;
mem[6263] = 80'h0010d845c0550102c000;
mem[6264] = 80'h00100001ffabffabffab;
mem[6265] = 80'h0010ffccf64307242f1b;
mem[6266] = 80'h0010c51aeeb33940e2b8;
mem[6267] = 80'h00104c84d563e1c60d95;
mem[6268] = 80'h01111200000000000000;
mem[6269] = 80'h00000000000000000000;
mem[6270] = 80'h10100000010000010010;
mem[6271] = 80'h00109400000208004500;
mem[6272] = 80'h0010002f61340000fffd;
mem[6273] = 80'h0010d844c0550102c000;
mem[6274] = 80'h00100001ffabffabffab;
mem[6275] = 80'h0010ffcbd287edf53b94;
mem[6276] = 80'h001045a201a2557c03c3;
mem[6277] = 80'h0010a915298990d04c96;
mem[6278] = 80'h01116500000000000000;
mem[6279] = 80'h00000000000000000000;
mem[6280] = 80'h00000000000000000000;
mem[6281] = 80'h00000000000000000000;
mem[6282] = 80'h10100000010000010010;
mem[6283] = 80'h00109400000208004500;
mem[6284] = 80'h0010002f61350000fffd;
mem[6285] = 80'h0010d843c0550102c000;
mem[6286] = 80'h00100001ffabffabffab;
mem[6287] = 80'h0010ffcaa359c12d4256;
mem[6288] = 80'h0010fa69d325b889d25a;
mem[6289] = 80'h0010f8f1a0f166337d98;
mem[6290] = 80'h0111c600000000000000;
mem[6291] = 80'h00000000000000000000;
mem[6292] = 80'h10100000010000010010;
mem[6293] = 80'h00109400000208004500;
mem[6294] = 80'h0010002f61360000fffd;
mem[6295] = 80'h0010d842c0550102c000;
mem[6296] = 80'h00100001ffabffabffab;
mem[6297] = 80'h0010ffc9313bb445c811;
mem[6298] = 80'h00103a35a4ad8e97a2d1;
mem[6299] = 80'h00100ab4bda3793b632b;
mem[6300] = 80'h01112900000000000000;
mem[6301] = 80'h00000000000000000000;
mem[6302] = 80'h00000000000000000000;
mem[6303] = 80'h00000000000000000000;
mem[6304] = 80'h00000000000000000000;
mem[6305] = 80'h10100000010000010010;
mem[6306] = 80'h00109400000208004500;
mem[6307] = 80'h0010002f61370000fffd;
mem[6308] = 80'h0010d841c0550102c000;
mem[6309] = 80'h00100001ffabffabffab;
mem[6310] = 80'h0010ffc840e5989db1d3;
mem[6311] = 80'h001085fe762a636272d8;
mem[6312] = 80'h00105b7feffd56559b38;
mem[6313] = 80'h01114c00000000000000;
mem[6314] = 80'h10100000010000010010;
mem[6315] = 80'h00109400000208004500;
mem[6316] = 80'h0010002f61380000fffd;
mem[6317] = 80'h0010d840c0550102c000;
mem[6318] = 80'h00100001ffabffabffab;
mem[6319] = 80'h0010ffc778b261e7e10e;
mem[6320] = 80'h00103b447a8f56ee6026;
mem[6321] = 80'h0010c197450fd09f3a4a;
mem[6322] = 80'h01117a00000000000000;
mem[6323] = 80'h00000000000000000000;
mem[6324] = 80'h00000000000000000000;
mem[6325] = 80'h00000000000000000000;
mem[6326] = 80'h10100000010000010010;
mem[6327] = 80'h00109400000208004500;
mem[6328] = 80'h0010002f61390000fffd;
mem[6329] = 80'h0010d83fc0550102c000;
mem[6330] = 80'h00100001ffabffabffab;
mem[6331] = 80'h0010ffc6096c4d3f98cc;
mem[6332] = 80'h0010848fa808bb1bb05f;
mem[6333] = 80'h001090544e59996b700f;
mem[6334] = 80'h01115d00000000000000;
mem[6335] = 80'h00000000000000000000;
mem[6336] = 80'h10100000010000010010;
mem[6337] = 80'h00109400000208004500;
mem[6338] = 80'h0010002f613a0000fffd;
mem[6339] = 80'h0010d83ec0550102c000;
mem[6340] = 80'h00100001ffabffabffab;
mem[6341] = 80'h0010ffc59b0e3857128b;
mem[6342] = 80'h001044d3df808d05c015;
mem[6343] = 80'h0010623436a60f950c35;
mem[6344] = 80'h01113e00000000000000;
mem[6345] = 80'h00000000000000000000;
mem[6346] = 80'h00000000000000000000;
mem[6347] = 80'h00000000000000000000;
mem[6348] = 80'h10100000010000010010;
mem[6349] = 80'h00109400000208004500;
mem[6350] = 80'h0010002f613b0000fffd;
mem[6351] = 80'h0010d83dc0550102c000;
mem[6352] = 80'h00100001ffabffabffab;
mem[6353] = 80'h0010ffc4ead0148f6b49;
mem[6354] = 80'h0010fb180d0760f0105c;
mem[6355] = 80'h001033f2a8333f1e4aa7;
mem[6356] = 80'h01119b00000000000000;
mem[6357] = 80'h00000000000000000000;
mem[6358] = 80'h00000000000000000000;
mem[6359] = 80'h00000000000000000000;
mem[6360] = 80'h10100000010000010010;
mem[6361] = 80'h00109400000208004500;
mem[6362] = 80'h0010002f613c0000fffd;
mem[6363] = 80'h0010d83cc0550102c000;
mem[6364] = 80'h00100001ffabffabffab;
mem[6365] = 80'h0010ffc3ce14fe5e7fc6;
mem[6366] = 80'h00107ba0e2160cccf167;
mem[6367] = 80'h0010d66e98a7e838e42a;
mem[6368] = 80'h01110700000000000000;
mem[6369] = 80'h00000000000000000000;
mem[6370] = 80'h10100000010000010010;
mem[6371] = 80'h00109400000208004500;
mem[6372] = 80'h0010002f613d0000fffd;
mem[6373] = 80'h0010d83bc0550102c000;
mem[6374] = 80'h00100001ffabffabffab;
mem[6375] = 80'h0010ffc2bfcad2860604;
mem[6376] = 80'h0010c46b3091e139213e;
mem[6377] = 80'h001087ab75c77256def4;
mem[6378] = 80'h01118200000000000000;
mem[6379] = 80'h00000000000000000000;
mem[6380] = 80'h10100000010000010010;
mem[6381] = 80'h00109400000208004500;
mem[6382] = 80'h0010002f613e0000fffd;
mem[6383] = 80'h0010d83ac0550102c000;
mem[6384] = 80'h00100001ffabffabffab;
mem[6385] = 80'h0010ffc12da8a7ee8c43;
mem[6386] = 80'h001004374719d7275275;
mem[6387] = 80'h001075a16cd5468592fc;
mem[6388] = 80'h0111d500000000000000;
mem[6389] = 80'h00000000000000000000;
mem[6390] = 80'h00000000000000000000;
mem[6391] = 80'h00000000000000000000;
mem[6392] = 80'h00000000000000000000;
mem[6393] = 80'h10100000010000010010;
mem[6394] = 80'h00109400000208004500;
mem[6395] = 80'h0010002f613f0000fffd;
mem[6396] = 80'h0010d839c0550102c000;
mem[6397] = 80'h00100001ffabffabffab;
mem[6398] = 80'h0010ffc05c768b36f581;
mem[6399] = 80'h0010bbfc959e3ad2823c;
mem[6400] = 80'h00102467f2fefc063d45;
mem[6401] = 80'h01110700000000000000;
mem[6402] = 80'h00000000000000000000;
mem[6403] = 80'h10100000010000010010;
mem[6404] = 80'h00109400000208004500;
mem[6405] = 80'h0010002f61400000fffd;
mem[6406] = 80'h0010d838c0550102c000;
mem[6407] = 80'h00100001ffabffabffab;
mem[6408] = 80'h0010ffbfcbd386ed1e21;
mem[6409] = 80'h0010715fcd20177b25b5;
mem[6410] = 80'h0010435a2653a9f377f9;
mem[6411] = 80'h0111b000000000000000;
mem[6412] = 80'h00000000000000000000;
mem[6413] = 80'h00000000000000000000;
mem[6414] = 80'h00000000000000000000;
mem[6415] = 80'h10100000010000010010;
mem[6416] = 80'h00109400000208004500;
mem[6417] = 80'h0010002f61410000fffd;
mem[6418] = 80'h0010d837c0550102c000;
mem[6419] = 80'h00100001ffabffabffab;
mem[6420] = 80'h0010ffbeba0daa3567e3;
mem[6421] = 80'h0010ce941fa7fa8ef5cc;
mem[6422] = 80'h001012992dea1476c1df;
mem[6423] = 80'h01113f00000000000000;
mem[6424] = 80'h00000000000000000000;
mem[6425] = 80'h10100000010000010010;
mem[6426] = 80'h00109400000208004500;
mem[6427] = 80'h0010002f61420000fffd;
mem[6428] = 80'h0010d836c0550102c000;
mem[6429] = 80'h00100001ffabffabffab;
mem[6430] = 80'h0010ffbd286fdf5deda4;
mem[6431] = 80'h00100ec8682fcc908547;
mem[6432] = 80'h0010e0dc3024304cf393;
mem[6433] = 80'h0111bc00000000000000;
mem[6434] = 80'h00000000000000000000;
mem[6435] = 80'h00000000000000000000;
mem[6436] = 80'h00000000000000000000;
mem[6437] = 80'h10100000010000010010;
mem[6438] = 80'h00109400000208004500;
mem[6439] = 80'h0010002f61430000fffd;
mem[6440] = 80'h0010d835c0550102c000;
mem[6441] = 80'h00100001ffabffabffab;
mem[6442] = 80'h0010ffbc59b1f3859466;
mem[6443] = 80'h0010b103baa8216555ce;
mem[6444] = 80'h0010b10cfab88fa400eb;
mem[6445] = 80'h0111ba00000000000000;
mem[6446] = 80'h00000000000000000000;
mem[6447] = 80'h10100000010000010010;
mem[6448] = 80'h00109400000208004500;
mem[6449] = 80'h0010002f61440000fffd;
mem[6450] = 80'h0010d834c0550102c000;
mem[6451] = 80'h00100001ffabffabffab;
mem[6452] = 80'h0010ffbb7d75195480e9;
mem[6453] = 80'h001031bb55b94d59b4b5;
mem[6454] = 80'h0010549d06710372b84d;
mem[6455] = 80'h0111b000000000000000;
mem[6456] = 80'h00000000000000000000;
mem[6457] = 80'h00000000000000000000;
mem[6458] = 80'h00000000000000000000;
mem[6459] = 80'h10100000010000010010;
mem[6460] = 80'h00109400000208004500;
mem[6461] = 80'h0010002f61450000fffd;
mem[6462] = 80'h0010d833c0550102c000;
mem[6463] = 80'h00100001ffabffabffab;
mem[6464] = 80'h0010ffba0cab358cf92b;
mem[6465] = 80'h00108e70873ea0ac64ac;
mem[6466] = 80'h0010055527857c606659;
mem[6467] = 80'h01119500000000000000;
mem[6468] = 80'h00000000000000000000;
mem[6469] = 80'h10100000010000010010;
mem[6470] = 80'h00109400000208004500;
mem[6471] = 80'h0010002f61460000fffd;
mem[6472] = 80'h0010d832c0550102c000;
mem[6473] = 80'h00100001ffabffabffab;
mem[6474] = 80'h0010ffb99ec940e4736c;
mem[6475] = 80'h00104e2cf0b696b21426;
mem[6476] = 80'h0010f7230b4cc0a6d2eb;
mem[6477] = 80'h0111ab00000000000000;
mem[6478] = 80'h00000000000000000000;
mem[6479] = 80'h00000000000000000000;
mem[6480] = 80'h00000000000000000000;
mem[6481] = 80'h10100000010000010010;
mem[6482] = 80'h00109400000208004500;
mem[6483] = 80'h0010002f61470000fffd;
mem[6484] = 80'h0010d831c0550102c000;
mem[6485] = 80'h00100001ffabffabffab;
mem[6486] = 80'h0010ffb8ef176c3c0aae;
mem[6487] = 80'h0010f1e722317b47c5af;
mem[6488] = 80'h0010a6c4f16fac6b3ef4;
mem[6489] = 80'h01113e00000000000000;
mem[6490] = 80'h00000000000000000000;
mem[6491] = 80'h10100000010000010010;
mem[6492] = 80'h00109400000208004500;
mem[6493] = 80'h0010002f61480000fffd;
mem[6494] = 80'h0010d830c0550102c000;
mem[6495] = 80'h00100001ffabffabffab;
mem[6496] = 80'h0010ffb7d74095465a73;
mem[6497] = 80'h00104f5d2e944ecbd751;
mem[6498] = 80'h00103c2c5b12fd525c2a;
mem[6499] = 80'h0111ac00000000000000;
mem[6500] = 80'h00000000000000000000;
mem[6501] = 80'h10100000010000010010;
mem[6502] = 80'h00109400000208004500;
mem[6503] = 80'h0010002f61490000fffd;
mem[6504] = 80'h0010d82fc0550102c000;
mem[6505] = 80'h00100001ffabffabffab;
mem[6506] = 80'h0010ffb6a69eb99e23b1;
mem[6507] = 80'h0010f096fc13a33e0728;
mem[6508] = 80'h00106def505a261a9c3b;
mem[6509] = 80'h01116b00000000000000;
mem[6510] = 80'h00000000000000000000;
mem[6511] = 80'h00000000000000000000;
mem[6512] = 80'h00000000000000000000;
mem[6513] = 80'h10100000010000010010;
mem[6514] = 80'h00109400000208004500;
mem[6515] = 80'h0010002f614a0000fffd;
mem[6516] = 80'h0010d82ec0550102c000;
mem[6517] = 80'h00100001ffabffabffab;
mem[6518] = 80'h0010ffb534fcccf6a9f6;
mem[6519] = 80'h001030ca8b9b952077e3;
mem[6520] = 80'h00109fa7814f69b1b75c;
mem[6521] = 80'h01113500000000000000;
mem[6522] = 80'h00000000000000000000;
mem[6523] = 80'h00000000000000000000;
mem[6524] = 80'h00000000000000000000;
mem[6525] = 80'h10100000010000010010;
mem[6526] = 80'h00109400000208004500;
mem[6527] = 80'h0010002f614b0000fffd;
mem[6528] = 80'h0010d82dc0550102c000;
mem[6529] = 80'h00100001ffabffabffab;
mem[6530] = 80'h0010ffb44522e02ed034;
mem[6531] = 80'h00108f01591c78d5a7aa;
mem[6532] = 80'h0010ce611fc613e904b0;
mem[6533] = 80'h0111e000000000000000;
mem[6534] = 80'h10100000010000010010;
mem[6535] = 80'h00109400000208004500;
mem[6536] = 80'h0010002f614c0000fffd;
mem[6537] = 80'h0010d82cc0550102c000;
mem[6538] = 80'h00100001ffabffabffab;
mem[6539] = 80'h0010ffb361e60affc4bb;
mem[6540] = 80'h00100fb9b60d14e94616;
mem[6541] = 80'h00102b7f206661b21312;
mem[6542] = 80'h01112e00000000000000;
mem[6543] = 80'h00000000000000000000;
mem[6544] = 80'h00000000000000000000;
mem[6545] = 80'h00000000000000000000;
mem[6546] = 80'h10100000010000010010;
mem[6547] = 80'h00109400000208004500;
mem[6548] = 80'h0010002f614d0000fffd;
mem[6549] = 80'h0010d82bc0550102c000;
mem[6550] = 80'h00100001ffabffabffab;
mem[6551] = 80'h0010ffb210382627bd79;
mem[6552] = 80'h0010b072648af91c9657;
mem[6553] = 80'h00107a3017d2d5474231;
mem[6554] = 80'h01117f00000000000000;
mem[6555] = 80'h00000000000000000000;
mem[6556] = 80'h10100000010000010010;
mem[6557] = 80'h00109400000208004500;
mem[6558] = 80'h0010002f614e0000fffd;
mem[6559] = 80'h0010d82ac0550102c000;
mem[6560] = 80'h00100001ffabffabffab;
mem[6561] = 80'h0010ffb1825a534f373e;
mem[6562] = 80'h0010702e1302cf02e684;
mem[6563] = 80'h001088f21cbc14b901e2;
mem[6564] = 80'h01110a00000000000000;
mem[6565] = 80'h00000000000000000000;
mem[6566] = 80'h00000000000000000000;
mem[6567] = 80'h00000000000000000000;
mem[6568] = 80'h10100000010000010010;
mem[6569] = 80'h00109400000208004500;
mem[6570] = 80'h0010002f614f0000fffd;
mem[6571] = 80'h0010d829c0550102c000;
mem[6572] = 80'h00100001ffabffabffab;
mem[6573] = 80'h0010ffb0f3847f974efc;
mem[6574] = 80'h0010cfe5c18522f736c5;
mem[6575] = 80'h0010d9bd2b514d037053;
mem[6576] = 80'h0111d600000000000000;
mem[6577] = 80'h00000000000000000000;
mem[6578] = 80'h10100000010000010010;
mem[6579] = 80'h00109400000208004500;
mem[6580] = 80'h0010002f61500000fffd;
mem[6581] = 80'h0010d828c0550102c000;
mem[6582] = 80'h00100001ffabffabffab;
mem[6583] = 80'h0010ffaff2f5a1bb9685;
mem[6584] = 80'h00100d5a0a48a41accf9;
mem[6585] = 80'h0010bc04c05dcfe48875;
mem[6586] = 80'h01115e00000000000000;
mem[6587] = 80'h00000000000000000000;
mem[6588] = 80'h00000000000000000000;
mem[6589] = 80'h00000000000000000000;
mem[6590] = 80'h00000000000000000000;
mem[6591] = 80'h10100000010000010010;
mem[6592] = 80'h00109400000208004500;
mem[6593] = 80'h0010002f61510000fffd;
mem[6594] = 80'h0010d827c0550102c000;
mem[6595] = 80'h00100001ffabffabffab;
mem[6596] = 80'h0010ffae832b8d63ef47;
mem[6597] = 80'h0010b291d8cf49ef1cb8;
mem[6598] = 80'h0010ed4bf72529a5c0dc;
mem[6599] = 80'h01119d00000000000000;
mem[6600] = 80'h10100000010000010010;
mem[6601] = 80'h00109400000208004500;
mem[6602] = 80'h0010002f61520000fffd;
mem[6603] = 80'h0010d826c0550102c000;
mem[6604] = 80'h00100001ffabffabffab;
mem[6605] = 80'h0010ffad1149f80b6500;
mem[6606] = 80'h001072cdaf477ff16c0b;
mem[6607] = 80'h00101f82d6688d802a51;
mem[6608] = 80'h01118100000000000000;
mem[6609] = 80'h00000000000000000000;
mem[6610] = 80'h00000000000000000000;
mem[6611] = 80'h00000000000000000000;
mem[6612] = 80'h10100000010000010010;
mem[6613] = 80'h00109400000208004500;
mem[6614] = 80'h0010002f61530000fffd;
mem[6615] = 80'h0010d825c0550102c000;
mem[6616] = 80'h00100001ffabffabffab;
mem[6617] = 80'h0010ffac6097d4d31cc2;
mem[6618] = 80'h0010cd067dc09204bc0b;
mem[6619] = 80'h00104ef31c5ba9f20803;
mem[6620] = 80'h01110500000000000000;
mem[6621] = 80'h00000000000000000000;
mem[6622] = 80'h10100000010000010010;
mem[6623] = 80'h00109400000208004500;
mem[6624] = 80'h0010002f61540000fffd;
mem[6625] = 80'h0010d824c0550102c000;
mem[6626] = 80'h00100001ffabffabffab;
mem[6627] = 80'h0010ffab44533e02084d;
mem[6628] = 80'h00104dbe92d1fe385d78;
mem[6629] = 80'h0010abeb498543eced5c;
mem[6630] = 80'h01110400000000000000;
mem[6631] = 80'h00000000000000000000;
mem[6632] = 80'h00000000000000000000;
mem[6633] = 80'h00000000000000000000;
mem[6634] = 80'h10100000010000010010;
mem[6635] = 80'h00109400000208004500;
mem[6636] = 80'h0010002f61550000fffd;
mem[6637] = 80'h0010d823c0550102c000;
mem[6638] = 80'h00100001ffabffabffab;
mem[6639] = 80'h0010ffaa358d12da718f;
mem[6640] = 80'h0010f275405613cd8df9;
mem[6641] = 80'h0010fab22a194c2ce8be;
mem[6642] = 80'h01115b00000000000000;
mem[6643] = 80'h00000000000000000000;
mem[6644] = 80'h10100000010000010010;
mem[6645] = 80'h00109400000208004500;
mem[6646] = 80'h0010002f61560000fffd;
mem[6647] = 80'h0010d822c0550102c000;
mem[6648] = 80'h00100001ffabffabffab;
mem[6649] = 80'h0010ffa9a7ef67b2fbc8;
mem[6650] = 80'h0010322937de25d3fd6a;
mem[6651] = 80'h0010087ded2871ebe9c2;
mem[6652] = 80'h0111c200000000000000;
mem[6653] = 80'h00000000000000000000;
mem[6654] = 80'h00000000000000000000;
mem[6655] = 80'h00000000000000000000;
mem[6656] = 80'h00000000000000000000;
mem[6657] = 80'h10100000010000010010;
mem[6658] = 80'h00109400000208004500;
mem[6659] = 80'h0010002f61570000fffd;
mem[6660] = 80'h0010d821c0550102c000;
mem[6661] = 80'h00100001ffabffabffab;
mem[6662] = 80'h0010ffa8d6314b6a820a;
mem[6663] = 80'h00108de2e559c8262d6b;
mem[6664] = 80'h0010593f16a383859357;
mem[6665] = 80'h01110900000000000000;
mem[6666] = 80'h10100000010000010010;
mem[6667] = 80'h00109400000208004500;
mem[6668] = 80'h0010002f61580000fffd;
mem[6669] = 80'h0010d820c0550102c000;
mem[6670] = 80'h00100001ffabffabffab;
mem[6671] = 80'h0010ffa7ee66b210d2d7;
mem[6672] = 80'h00103358e9fcfdaa3f9d;
mem[6673] = 80'h0010c35e150d59fb205d;
mem[6674] = 80'h0111e100000000000000;
mem[6675] = 80'h00000000000000000000;
mem[6676] = 80'h00000000000000000000;
mem[6677] = 80'h00000000000000000000;
mem[6678] = 80'h10100000010000010010;
mem[6679] = 80'h00109400000208004500;
mem[6680] = 80'h0010002f61590000fffd;
mem[6681] = 80'h0010d81fc0550102c000;
mem[6682] = 80'h00100001ffabffabffab;
mem[6683] = 80'h0010ffa69fb89ec8ab15;
mem[6684] = 80'h00108c933b7b105fee1f;
mem[6685] = 80'h0010926515cfa70bb572;
mem[6686] = 80'h01112300000000000000;
mem[6687] = 80'h00000000000000000000;
mem[6688] = 80'h10100000010000010010;
mem[6689] = 80'h00109400000208004500;
mem[6690] = 80'h0010002f615a0000fffd;
mem[6691] = 80'h0010d81ec0550102c000;
mem[6692] = 80'h00100001ffabffabffab;
mem[6693] = 80'h0010ffa50ddaeba02152;
mem[6694] = 80'h00104ccf4cf326419eac;
mem[6695] = 80'h001060ac3430f12400bf;
mem[6696] = 80'h0111ba00000000000000;
mem[6697] = 80'h00000000000000000000;
mem[6698] = 80'h00000000000000000000;
mem[6699] = 80'h00000000000000000000;
mem[6700] = 80'h10100000010000010010;
mem[6701] = 80'h00109400000208004500;
mem[6702] = 80'h0010002f615b0000fffd;
mem[6703] = 80'h0010d81dc0550102c000;
mem[6704] = 80'h00100001ffabffabffab;
mem[6705] = 80'h0010ffa47c04c7785890;
mem[6706] = 80'h0010f3049e74cbb44eed;
mem[6707] = 80'h001031e3034f82d050c2;
mem[6708] = 80'h0111fe00000000000000;
mem[6709] = 80'h00000000000000000000;
mem[6710] = 80'h00000000000000000000;
mem[6711] = 80'h00000000000000000000;
mem[6712] = 80'h10100000010000010010;
mem[6713] = 80'h00109400000208004500;
mem[6714] = 80'h0010002f615c0000fffd;
mem[6715] = 80'h0010d81cc0550102c000;
mem[6716] = 80'h00100001ffabffabffab;
mem[6717] = 80'h0010ffa358c02da94c1f;
mem[6718] = 80'h001073bc7165a788afde;
mem[6719] = 80'h0010d4f69a53814be700;
mem[6720] = 80'h0111ba00000000000000;
mem[6721] = 80'h00000000000000000000;
mem[6722] = 80'h10100000010000010010;
mem[6723] = 80'h00109400000208004500;
mem[6724] = 80'h0010002f615d0000fffd;
mem[6725] = 80'h0010d81bc0550102c000;
mem[6726] = 80'h00100001ffabffabffab;
mem[6727] = 80'h0010ffa2291e017135dd;
mem[6728] = 80'h0010cc77a3e24a7d7f9f;
mem[6729] = 80'h001085b9adc031c2c08b;
mem[6730] = 80'h01113600000000000000;
mem[6731] = 80'h00000000000000000000;
mem[6732] = 80'h10100000010000010010;
mem[6733] = 80'h00109400000208004500;
mem[6734] = 80'h0010002f615e0000fffd;
mem[6735] = 80'h0010d81ac0550102c000;
mem[6736] = 80'h00100001ffabffabffab;
mem[6737] = 80'h0010ffa1bb7c7419bf9a;
mem[6738] = 80'h00100c2bd46a7c630fcc;
mem[6739] = 80'h001077603e07eef1943a;
mem[6740] = 80'h0111ac00000000000000;
mem[6741] = 80'h00000000000000000000;
mem[6742] = 80'h00000000000000000000;
mem[6743] = 80'h00000000000000000000;
mem[6744] = 80'h00000000000000000000;
mem[6745] = 80'h10100000010000010010;
mem[6746] = 80'h00109400000208004500;
mem[6747] = 80'h0010002f615f0000fffd;
mem[6748] = 80'h0010d819c0550102c000;
mem[6749] = 80'h00100001ffabffabffab;
mem[6750] = 80'h0010ffa0caa258c1c658;
mem[6751] = 80'h0010b3e006ed9196df8c;
mem[6752] = 80'h0010261c38958bb8f728;
mem[6753] = 80'h0111fb00000000000000;
mem[6754] = 80'h00000000000000000000;
mem[6755] = 80'h10100000010000010010;
mem[6756] = 80'h00109400000208004500;
mem[6757] = 80'h0010002f61600000fffd;
mem[6758] = 80'h0010d818c0550102c000;
mem[6759] = 80'h00100001ffabffabffab;
mem[6760] = 80'h0010ff9fb99fc8400f69;
mem[6761] = 80'h0010895443f171b8e425;
mem[6762] = 80'h0010bd4741ab4ca352fa;
mem[6763] = 80'h0111f200000000000000;
mem[6764] = 80'h00000000000000000000;
mem[6765] = 80'h00000000000000000000;
mem[6766] = 80'h00000000000000000000;
mem[6767] = 80'h10100000010000010010;
mem[6768] = 80'h00109400000208004500;
mem[6769] = 80'h0010002f61610000fffd;
mem[6770] = 80'h0010d817c0550102c000;
mem[6771] = 80'h00100001ffabffabffab;
mem[6772] = 80'h0010ff9ec841e49876ab;
mem[6773] = 80'h0010369f91769c4d3464;
mem[6774] = 80'h0010ec08760ae1acfca7;
mem[6775] = 80'h01118000000000000000;
mem[6776] = 80'h00000000000000000000;
mem[6777] = 80'h10100000010000010010;
mem[6778] = 80'h00109400000208004500;
mem[6779] = 80'h0010002f61620000fffd;
mem[6780] = 80'h0010d816c0550102c000;
mem[6781] = 80'h00100001ffabffabffab;
mem[6782] = 80'h0010ff9d5a2391f0fcec;
mem[6783] = 80'h0010f6c3e6feaa5344d7;
mem[6784] = 80'h00101ec157b2d300358d;
mem[6785] = 80'h0111ec00000000000000;
mem[6786] = 80'h00000000000000000000;
mem[6787] = 80'h00000000000000000000;
mem[6788] = 80'h00000000000000000000;
mem[6789] = 80'h10100000010000010010;
mem[6790] = 80'h00109400000208004500;
mem[6791] = 80'h0010002f61630000fffd;
mem[6792] = 80'h0010d815c0550102c000;
mem[6793] = 80'h00100001ffabffabffab;
mem[6794] = 80'h0010ff9c2bfdbd28852e;
mem[6795] = 80'h00104908347947a69756;
mem[6796] = 80'h00104fc164cf8020c3d6;
mem[6797] = 80'h01114500000000000000;
mem[6798] = 80'h00000000000000000000;
mem[6799] = 80'h10100000010000010010;
mem[6800] = 80'h00109400000208004500;
mem[6801] = 80'h0010002f61640000fffd;
mem[6802] = 80'h0010d814c0550102c000;
mem[6803] = 80'h00100001ffabffabffab;
mem[6804] = 80'h0010ff9b0f3957f991a1;
mem[6805] = 80'h0010c9b0db682b9a7625;
mem[6806] = 80'h0010aad931dde3f885a2;
mem[6807] = 80'h0111b700000000000000;
mem[6808] = 80'h00000000000000000000;
mem[6809] = 80'h00000000000000000000;
mem[6810] = 80'h00000000000000000000;
mem[6811] = 80'h10100000010000010010;
mem[6812] = 80'h00109400000208004500;
mem[6813] = 80'h0010002f61650000fffd;
mem[6814] = 80'h0010d813c0550102c000;
mem[6815] = 80'h00100001ffabffabffab;
mem[6816] = 80'h0010ff9a7ee77b21e863;
mem[6817] = 80'h0010767b09efc66fa623;
mem[6818] = 80'h0010fb025df7d7cf7d6d;
mem[6819] = 80'h0111a400000000000000;
mem[6820] = 80'h00000000000000000000;
mem[6821] = 80'h10100000010000010010;
mem[6822] = 80'h00109400000208004500;
mem[6823] = 80'h0010002f61660000fffd;
mem[6824] = 80'h0010d812c0550102c000;
mem[6825] = 80'h00100001ffabffabffab;
mem[6826] = 80'h0010ff99ec850e496224;
mem[6827] = 80'h0010b6277e67f071d6a8;
mem[6828] = 80'h0010094740825d69b67e;
mem[6829] = 80'h01111100000000000000;
mem[6830] = 80'h00000000000000000000;
mem[6831] = 80'h00000000000000000000;
mem[6832] = 80'h00000000000000000000;
mem[6833] = 80'h10100000010000010010;
mem[6834] = 80'h00109400000208004500;
mem[6835] = 80'h0010002f61670000fffd;
mem[6836] = 80'h0010d811c0550102c000;
mem[6837] = 80'h00100001ffabffabffab;
mem[6838] = 80'h0010ff989d5b22911be6;
mem[6839] = 80'h001009ecace01d840631;
mem[6840] = 80'h00105894f97df772e2df;
mem[6841] = 80'h01117300000000000000;
mem[6842] = 80'h00000000000000000000;
mem[6843] = 80'h10100000010000010010;
mem[6844] = 80'h00109400000208004500;
mem[6845] = 80'h0010002f61680000fffd;
mem[6846] = 80'h0010d810c0550102c000;
mem[6847] = 80'h00100001ffabffabffab;
mem[6848] = 80'h0010ff97a50cdbeb4b3b;
mem[6849] = 80'h0010b756a045280814cf;
mem[6850] = 80'h0010c27c5344891337c5;
mem[6851] = 80'h0111de00000000000000;
mem[6852] = 80'h00000000000000000000;
mem[6853] = 80'h10100000010000010010;
mem[6854] = 80'h00109400000208004500;
mem[6855] = 80'h0010002f61690000fffd;
mem[6856] = 80'h0010d80fc0550102c000;
mem[6857] = 80'h00100001ffabffabffab;
mem[6858] = 80'h0010ff96d4d2f73332f9;
mem[6859] = 80'h0010089d72c2c5fdc4c6;
mem[6860] = 80'h001093b7018e658c9827;
mem[6861] = 80'h01110500000000000000;
mem[6862] = 80'h00000000000000000000;
mem[6863] = 80'h00000000000000000000;
mem[6864] = 80'h00000000000000000000;
mem[6865] = 80'h10100000010000010010;
mem[6866] = 80'h00109400000208004500;
mem[6867] = 80'h0010002f616a0000fffd;
mem[6868] = 80'h0010d80ec0550102c000;
mem[6869] = 80'h00100001ffabffabffab;
mem[6870] = 80'h0010ff9546b0825bb8be;
mem[6871] = 80'h0010c8c1054af3e3b44d;
mem[6872] = 80'h001061f21c7089c7d692;
mem[6873] = 80'h0111cc00000000000000;
mem[6874] = 80'h00000000000000000000;
mem[6875] = 80'h00000000000000000000;
mem[6876] = 80'h00000000000000000000;
mem[6877] = 80'h10100000010000010010;
mem[6878] = 80'h00109400000208004500;
mem[6879] = 80'h0010002f616b0000fffd;
mem[6880] = 80'h0010d80dc0550102c000;
mem[6881] = 80'h00100001ffabffabffab;
mem[6882] = 80'h0010ff94376eae83c17c;
mem[6883] = 80'h0010770ad7cd1e166434;
mem[6884] = 80'h0010303117a93fd43b6b;
mem[6885] = 80'h0111f900000000000000;
mem[6886] = 80'h10100000010000010010;
mem[6887] = 80'h00109400000208004500;
mem[6888] = 80'h0010002f616c0000fffd;
mem[6889] = 80'h0010d80cc0550102c000;
mem[6890] = 80'h00100001ffabffabffab;
mem[6891] = 80'h0010ff9313aa4452d5f3;
mem[6892] = 80'h0010f7b238dc722a848e;
mem[6893] = 80'h0010d5b2be811622a3b0;
mem[6894] = 80'h0111fe00000000000000;
mem[6895] = 80'h00000000000000000000;
mem[6896] = 80'h00000000000000000000;
mem[6897] = 80'h00000000000000000000;
mem[6898] = 80'h10100000010000010010;
mem[6899] = 80'h00109400000208004500;
mem[6900] = 80'h0010002f616d0000fffd;
mem[6901] = 80'h0010d80bc0550102c000;
mem[6902] = 80'h00100001ffabffabffab;
mem[6903] = 80'h0010ff926274688aac31;
mem[6904] = 80'h00104879ea5b9fdf54c7;
mem[6905] = 80'h00108474204cbc3810ca;
mem[6906] = 80'h01110100000000000000;
mem[6907] = 80'h00000000000000000000;
mem[6908] = 80'h10100000010000010010;
mem[6909] = 80'h00109400000208004500;
mem[6910] = 80'h0010002f616e0000fffd;
mem[6911] = 80'h0010d80ac0550102c000;
mem[6912] = 80'h00100001ffabffabffab;
mem[6913] = 80'h0010ff91f0161de22676;
mem[6914] = 80'h001088259dd3a9c1240c;
mem[6915] = 80'h0010763cf1fb6f973a25;
mem[6916] = 80'h01113a00000000000000;
mem[6917] = 80'h00000000000000000000;
mem[6918] = 80'h00000000000000000000;
mem[6919] = 80'h00000000000000000000;
mem[6920] = 80'h10100000010000010010;
mem[6921] = 80'h00109400000208004500;
mem[6922] = 80'h0010002f616f0000fffd;
mem[6923] = 80'h0010d809c0550102c000;
mem[6924] = 80'h00100001ffabffabffab;
mem[6925] = 80'h0010ff9081c8313a5fb4;
mem[6926] = 80'h001037ee4f544434f455;
mem[6927] = 80'h001027f91cf2e859e492;
mem[6928] = 80'h01115000000000000000;
mem[6929] = 80'h00000000000000000000;
mem[6930] = 80'h10100000010000010010;
mem[6931] = 80'h00109400000208004500;
mem[6932] = 80'h0010002f61700000fffd;
mem[6933] = 80'h0010d808c0550102c000;
mem[6934] = 80'h00100001ffabffabffab;
mem[6935] = 80'h0010ff8f80b9ef1687cd;
mem[6936] = 80'h0010f5518499c2d90161;
mem[6937] = 80'h001042e56fc7177e6e2a;
mem[6938] = 80'h01116b00000000000000;
mem[6939] = 80'h00000000000000000000;
mem[6940] = 80'h00000000000000000000;
mem[6941] = 80'h00000000000000000000;
mem[6942] = 80'h00000000000000000000;
mem[6943] = 80'h10100000010000010010;
mem[6944] = 80'h00109400000208004500;
mem[6945] = 80'h0010002f61710000fffd;
mem[6946] = 80'h0010d807c0550102c000;
mem[6947] = 80'h00100001ffabffabffab;
mem[6948] = 80'h0010ff8ef167c3cefe0f;
mem[6949] = 80'h00104a9a561e2f2cd128;
mem[6950] = 80'h00101323f1f9a6d81704;
mem[6951] = 80'h01115100000000000000;
mem[6952] = 80'h10100000010000010010;
mem[6953] = 80'h00109400000208004500;
mem[6954] = 80'h0010002f61720000fffd;
mem[6955] = 80'h0010d806c0550102c000;
mem[6956] = 80'h00100001ffabffabffab;
mem[6957] = 80'h0010ff8d6305b6a67448;
mem[6958] = 80'h00108ac621961932a1e0;
mem[6959] = 80'h0010e13e73cfb51a4baa;
mem[6960] = 80'h0111c700000000000000;
mem[6961] = 80'h00000000000000000000;
mem[6962] = 80'h00000000000000000000;
mem[6963] = 80'h00000000000000000000;
mem[6964] = 80'h10100000010000010010;
mem[6965] = 80'h00109400000208004500;
mem[6966] = 80'h0010002f61730000fffd;
mem[6967] = 80'h0010d805c0550102c000;
mem[6968] = 80'h00100001ffabffabffab;
mem[6969] = 80'h0010ff8c12db9a7e0d8a;
mem[6970] = 80'h0010350df311f4c77199;
mem[6971] = 80'h0010b0fd78118de99e12;
mem[6972] = 80'h0111b700000000000000;
mem[6973] = 80'h00000000000000000000;
mem[6974] = 80'h10100000010000010010;
mem[6975] = 80'h00109400000208004500;
mem[6976] = 80'h0010002f61740000fffd;
mem[6977] = 80'h0010d804c0550102c000;
mem[6978] = 80'h00100001ffabffabffab;
mem[6979] = 80'h0010ff8b361f70af1905;
mem[6980] = 80'h0010b5b51c0098fb90e2;
mem[6981] = 80'h0010556c84a06a116d32;
mem[6982] = 80'h01118000000000000000;
mem[6983] = 80'h00000000000000000000;
mem[6984] = 80'h00000000000000000000;
mem[6985] = 80'h00000000000000000000;
mem[6986] = 80'h10100000010000010010;
mem[6987] = 80'h00109400000208004500;
mem[6988] = 80'h0010002f61750000fffd;
mem[6989] = 80'h0010d803c0550102c000;
mem[6990] = 80'h00100001ffabffabffab;
mem[6991] = 80'h0010ff8a47c15c7760c7;
mem[6992] = 80'h00100a7ece87750e476b;
mem[6993] = 80'h00100439debc82055aa5;
mem[6994] = 80'h01119200000000000000;
mem[6995] = 80'h00000000000000000000;
mem[6996] = 80'h10100000010000010010;
mem[6997] = 80'h00109400000208004500;
mem[6998] = 80'h0010002f61760000fffd;
mem[6999] = 80'h0010d802c0550102c000;
mem[7000] = 80'h00100001ffabffabffab;
mem[7001] = 80'h0010ff89d5a3291fea80;
mem[7002] = 80'h0010ca22b90f431037e0;
mem[7003] = 80'h0010f67cc3925efde1f1;
mem[7004] = 80'h0111fc00000000000000;
mem[7005] = 80'h00000000000000000000;
mem[7006] = 80'h00000000000000000000;
mem[7007] = 80'h00000000000000000000;
mem[7008] = 80'h00000000000000000000;
mem[7009] = 80'h10100000010000010010;
mem[7010] = 80'h00109400000208004500;
mem[7011] = 80'h0010002f61770000fffd;
mem[7012] = 80'h0010d801c0550102c000;
mem[7013] = 80'h00100001ffabffabffab;
mem[7014] = 80'h0010ff88a47d05c79342;
mem[7015] = 80'h001075e96b88aee5e7f9;
mem[7016] = 80'h0010a7b4e2e9bfbf5d19;
mem[7017] = 80'h01114a00000000000000;
mem[7018] = 80'h10100000010000010010;
mem[7019] = 80'h00109400000208004500;
mem[7020] = 80'h0010002f61780000fffd;
mem[7021] = 80'h0010d800c0550102c000;
mem[7022] = 80'h00100001ffabffabffab;
mem[7023] = 80'h0010ff879c2afcbdc39f;
mem[7024] = 80'h0010cb53672d9b69f506;
mem[7025] = 80'h00103d6f798f2942a89a;
mem[7026] = 80'h01117800000000000000;
mem[7027] = 80'h00000000000000000000;
mem[7028] = 80'h00000000000000000000;
mem[7029] = 80'h00000000000000000000;
mem[7030] = 80'h10100000010000010010;
mem[7031] = 80'h00109400000208004500;
mem[7032] = 80'h0010002f61790000fffd;
mem[7033] = 80'h0010d7ffc0550102c000;
mem[7034] = 80'h00100001ffabffabffab;
mem[7035] = 80'h0010ff86edf4d065ba5d;
mem[7036] = 80'h00107498b5aa769c258f;
mem[7037] = 80'h00106cbfb392a092643e;
mem[7038] = 80'h01119f00000000000000;
mem[7039] = 80'h00000000000000000000;
mem[7040] = 80'h10100000010000010010;
mem[7041] = 80'h00109400000208004500;
mem[7042] = 80'h0010002f617a0000fffd;
mem[7043] = 80'h0010d7fec0550102c000;
mem[7044] = 80'h00100001ffabffabffab;
mem[7045] = 80'h0010ff857f96a50d301a;
mem[7046] = 80'h0010b4c4c22240825504;
mem[7047] = 80'h00109efaae53513c6c53;
mem[7048] = 80'h01116d00000000000000;
mem[7049] = 80'h00000000000000000000;
mem[7050] = 80'h00000000000000000000;
mem[7051] = 80'h00000000000000000000;
mem[7052] = 80'h10100000010000010010;
mem[7053] = 80'h00109400000208004500;
mem[7054] = 80'h0010002f617b0000fffd;
mem[7055] = 80'h0010d7fdc0550102c000;
mem[7056] = 80'h00100001ffabffabffab;
mem[7057] = 80'h0010ff840e4889d549d8;
mem[7058] = 80'h00100b0f10a5ad77857d;
mem[7059] = 80'h0010cf39a5a25ab4e027;
mem[7060] = 80'h0111b000000000000000;
mem[7061] = 80'h00000000000000000000;
mem[7062] = 80'h00000000000000000000;
mem[7063] = 80'h00000000000000000000;
mem[7064] = 80'h10100000010000010010;
mem[7065] = 80'h00109400000208004500;
mem[7066] = 80'h0010002f617c0000fffd;
mem[7067] = 80'h0010d7fcc0550102c000;
mem[7068] = 80'h00100001ffabffabffab;
mem[7069] = 80'h0010ff832a8c63045d57;
mem[7070] = 80'h00108bb7ffb4c14b6446;
mem[7071] = 80'h00102aa595f0a39533dc;
mem[7072] = 80'h01116d00000000000000;
mem[7073] = 80'h00000000000000000000;
mem[7074] = 80'h10100000010000010010;
mem[7075] = 80'h00109400000208004500;
mem[7076] = 80'h0010002f617d0000fffd;
mem[7077] = 80'h0010d7fbc0550102c000;
mem[7078] = 80'h00100001ffabffabffab;
mem[7079] = 80'h0010ff825b524fdc2495;
mem[7080] = 80'h0010347c2d332cbeb40f;
mem[7081] = 80'h00107b630bd966aecab9;
mem[7082] = 80'h01117500000000000000;
mem[7083] = 80'h00000000000000000000;
mem[7084] = 80'h10100000010000010010;
mem[7085] = 80'h00109400000208004500;
mem[7086] = 80'h0010002f617e0000fffd;
mem[7087] = 80'h0010d7fac0550102c000;
mem[7088] = 80'h00100001ffabffabffab;
mem[7089] = 80'h0010ff81c9303ab4aed2;
mem[7090] = 80'h0010f4205abb1aa0c543;
mem[7091] = 80'h0010899ee567afe391af;
mem[7092] = 80'h0111c200000000000000;
mem[7093] = 80'h00000000000000000000;
mem[7094] = 80'h00000000000000000000;
mem[7095] = 80'h00000000000000000000;
mem[7096] = 80'h00000000000000000000;
mem[7097] = 80'h10100000010000010010;
mem[7098] = 80'h00109400000208004500;
mem[7099] = 80'h0010002f617f0000fffd;
mem[7100] = 80'h0010d7f9c0550102c000;
mem[7101] = 80'h00100001ffabffabffab;
mem[7102] = 80'h0010ff80b8ee166cd710;
mem[7103] = 80'h00104beb883cf7551502;
mem[7104] = 80'h0010d8d1d2c1cdb39f98;
mem[7105] = 80'h0111bc00000000000000;
mem[7106] = 80'h00000000000000000000;
mem[7107] = 80'h10100000010000010010;
mem[7108] = 80'h00109400000208004500;
mem[7109] = 80'h0010002f61800000fffd;
mem[7110] = 80'h0010d7f8c0550102c000;
mem[7111] = 80'h00100001ffabffabffab;
mem[7112] = 80'h0010ff7f97a40ddb0051;
mem[7113] = 80'h0010dead3941ac065aa2;
mem[7114] = 80'h0010178794908f0876c5;
mem[7115] = 80'h01117000000000000000;
mem[7116] = 80'h00000000000000000000;
mem[7117] = 80'h00000000000000000000;
mem[7118] = 80'h00000000000000000000;
mem[7119] = 80'h10100000010000010010;
mem[7120] = 80'h00109400000208004500;
mem[7121] = 80'h0010002f61810000fffd;
mem[7122] = 80'h0010d7f7c0550102c000;
mem[7123] = 80'h00100001ffabffabffab;
mem[7124] = 80'h0010ff7ee67a21037993;
mem[7125] = 80'h00106166ebc641f38ae3;
mem[7126] = 80'h001046c8a3a37a59e95f;
mem[7127] = 80'h01112400000000000000;
mem[7128] = 80'h00000000000000000000;
mem[7129] = 80'h10100000010000010010;
mem[7130] = 80'h00109400000208004500;
mem[7131] = 80'h0010002f61820000fffd;
mem[7132] = 80'h0010d7f6c0550102c000;
mem[7133] = 80'h00100001ffabffabffab;
mem[7134] = 80'h0010ff7d7418546bf3d4;
mem[7135] = 80'h0010a13a9c4e77edfaa0;
mem[7136] = 80'h0010b41243ff9b6c88ee;
mem[7137] = 80'h0111aa00000000000000;
mem[7138] = 80'h00000000000000000000;
mem[7139] = 80'h00000000000000000000;
mem[7140] = 80'h00000000000000000000;
mem[7141] = 80'h10100000010000010010;
mem[7142] = 80'h00109400000208004500;
mem[7143] = 80'h0010002f61830000fffd;
mem[7144] = 80'h0010d7f5c0550102c000;
mem[7145] = 80'h00100001ffabffabffab;
mem[7146] = 80'h0010ff7c05c678b38a16;
mem[7147] = 80'h00101ef14ec99a182ae1;
mem[7148] = 80'h0010e55d74e16a7260c3;
mem[7149] = 80'h01119100000000000000;
mem[7150] = 80'h00000000000000000000;
mem[7151] = 80'h10100000010000010010;
mem[7152] = 80'h00109400000208004500;
mem[7153] = 80'h0010002f61840000fffd;
mem[7154] = 80'h0010d7f4c0550102c000;
mem[7155] = 80'h00100001ffabffabffab;
mem[7156] = 80'h0010ff7b210292629e99;
mem[7157] = 80'h00109e49a1d8f624cba2;
mem[7158] = 80'h00100040b45bf7d44210;
mem[7159] = 80'h01119700000000000000;
mem[7160] = 80'h00000000000000000000;
mem[7161] = 80'h00000000000000000000;
mem[7162] = 80'h00000000000000000000;
mem[7163] = 80'h10100000010000010010;
mem[7164] = 80'h00109400000208004500;
mem[7165] = 80'h0010002f61850000fffd;
mem[7166] = 80'h0010d7f3c0550102c000;
mem[7167] = 80'h00100001ffabffabffab;
mem[7168] = 80'h0010ff7a50dcbebae75b;
mem[7169] = 80'h00102182735f1bd11ba2;
mem[7170] = 80'h001051317e0c6d19085a;
mem[7171] = 80'h01110600000000000000;
mem[7172] = 80'h00000000000000000000;
mem[7173] = 80'h10100000010000010010;
mem[7174] = 80'h00109400000208004500;
mem[7175] = 80'h0010002f61860000fffd;
mem[7176] = 80'h0010d7f2c0550102c000;
mem[7177] = 80'h00100001ffabffabffab;
mem[7178] = 80'h0010ff79c2becbd26d1c;
mem[7179] = 80'h0010e1de04d72dcf6b21;
mem[7180] = 80'h0010a3fdca34164e2d8f;
mem[7181] = 80'h01119600000000000000;
mem[7182] = 80'h00000000000000000000;
mem[7183] = 80'h00000000000000000000;
mem[7184] = 80'h00000000000000000000;
mem[7185] = 80'h10100000010000010010;
mem[7186] = 80'h00109400000208004500;
mem[7187] = 80'h0010002f61870000fffd;
mem[7188] = 80'h0010d7f1c0550102c000;
mem[7189] = 80'h00100001ffabffabffab;
mem[7190] = 80'h0010ff78b360e70a14de;
mem[7191] = 80'h00105e15d650c03ab8a0;
mem[7192] = 80'h0010f2fdf9fdb67413c9;
mem[7193] = 80'h01119b00000000000000;
mem[7194] = 80'h00000000000000000000;
mem[7195] = 80'h10100000010000010010;
mem[7196] = 80'h00109400000208004500;
mem[7197] = 80'h0010002f61880000fffd;
mem[7198] = 80'h0010d7f0c0550102c000;
mem[7199] = 80'h00100001ffabffabffab;
mem[7200] = 80'h0010ff778b371e704403;
mem[7201] = 80'h0010e0afdaf5f5b6aa46;
mem[7202] = 80'h0010689f899ac4ab9c22;
mem[7203] = 80'h0111f600000000000000;
mem[7204] = 80'h00000000000000000000;
mem[7205] = 80'h10100000010000010010;
mem[7206] = 80'h00109400000208004500;
mem[7207] = 80'h0010002f61890000fffd;
mem[7208] = 80'h0010d7efc0550102c000;
mem[7209] = 80'h00100001ffabffabffab;
mem[7210] = 80'h0010ff76fae932a83dc1;
mem[7211] = 80'h00105f64087218437a47;
mem[7212] = 80'h001039dd72f7ed163223;
mem[7213] = 80'h01118d00000000000000;
mem[7214] = 80'h00000000000000000000;
mem[7215] = 80'h00000000000000000000;
mem[7216] = 80'h00000000000000000000;
mem[7217] = 80'h10100000010000010010;
mem[7218] = 80'h00109400000208004500;
mem[7219] = 80'h0010002f618a0000fffd;
mem[7220] = 80'h0010d7eec0550102c000;
mem[7221] = 80'h00100001ffabffabffab;
mem[7222] = 80'h0010ff75688b47c0b786;
mem[7223] = 80'h00109f387ffa2e5d0ac4;
mem[7224] = 80'h0010cb11c651ae4b0836;
mem[7225] = 80'h0111da00000000000000;
mem[7226] = 80'h00000000000000000000;
mem[7227] = 80'h00000000000000000000;
mem[7228] = 80'h00000000000000000000;
mem[7229] = 80'h10100000010000010010;
mem[7230] = 80'h00109400000208004500;
mem[7231] = 80'h0010002f618b0000fffd;
mem[7232] = 80'h0010d7edc0550102c000;
mem[7233] = 80'h00100001ffabffabffab;
mem[7234] = 80'h0010ff7419556b18ce44;
mem[7235] = 80'h001020f3ad7dc3a8da46;
mem[7236] = 80'h00109a1df65ab0e47489;
mem[7237] = 80'h0111fd00000000000000;
mem[7238] = 80'h10100000010000010010;
mem[7239] = 80'h00109400000208004500;
mem[7240] = 80'h0010002f618c0000fffd;
mem[7241] = 80'h0010d7ecc0550102c000;
mem[7242] = 80'h00100001ffabffabffab;
mem[7243] = 80'h0010ff733d9181c9dacb;
mem[7244] = 80'h0010a04b426caf943b05;
mem[7245] = 80'h00107f003613e38b0b17;
mem[7246] = 80'h0111b800000000000000;
mem[7247] = 80'h00000000000000000000;
mem[7248] = 80'h00000000000000000000;
mem[7249] = 80'h00000000000000000000;
mem[7250] = 80'h10100000010000010010;
mem[7251] = 80'h00109400000208004500;
mem[7252] = 80'h0010002f618d0000fffd;
mem[7253] = 80'h0010d7ebc0550102c000;
mem[7254] = 80'h00100001ffabffabffab;
mem[7255] = 80'h0010ff724c4fad11a309;
mem[7256] = 80'h00101f8090eb4261eb44;
mem[7257] = 80'h00102e4f01c255b0a4b0;
mem[7258] = 80'h01111f00000000000000;
mem[7259] = 80'h00000000000000000000;
mem[7260] = 80'h10100000010000010010;
mem[7261] = 80'h00109400000208004500;
mem[7262] = 80'h0010002f618e0000fffd;
mem[7263] = 80'h0010d7eac0550102c000;
mem[7264] = 80'h00100001ffabffabffab;
mem[7265] = 80'h0010ff71de2dd879294e;
mem[7266] = 80'h0010dfdce763747f9b87;
mem[7267] = 80'h0010dc8e79c1f2b54d35;
mem[7268] = 80'h01115900000000000000;
mem[7269] = 80'h00000000000000000000;
mem[7270] = 80'h00000000000000000000;
mem[7271] = 80'h00000000000000000000;
mem[7272] = 80'h10100000010000010010;
mem[7273] = 80'h00109400000208004500;
mem[7274] = 80'h0010002f618f0000fffd;
mem[7275] = 80'h0010d7e9c0550102c000;
mem[7276] = 80'h00100001ffabffabffab;
mem[7277] = 80'h0010ff70aff3f4a1508c;
mem[7278] = 80'h0010601735e4998a4bc6;
mem[7279] = 80'h00108dc14e5fb36c8efa;
mem[7280] = 80'h01119200000000000000;
mem[7281] = 80'h00000000000000000000;
mem[7282] = 80'h10100000010000010010;
mem[7283] = 80'h00109400000208004500;
mem[7284] = 80'h0010002f61900000fffd;
mem[7285] = 80'h0010d7e8c0550102c000;
mem[7286] = 80'h00100001ffabffabffab;
mem[7287] = 80'h0010ff6fae822a8d88f5;
mem[7288] = 80'h0010a2a8fe291f67bfea;
mem[7289] = 80'h0010e860d7055e184a01;
mem[7290] = 80'h0111ba00000000000000;
mem[7291] = 80'h00000000000000000000;
mem[7292] = 80'h00000000000000000000;
mem[7293] = 80'h00000000000000000000;
mem[7294] = 80'h00000000000000000000;
mem[7295] = 80'h10100000010000010010;
mem[7296] = 80'h00109400000208004500;
mem[7297] = 80'h0010002f61910000fffd;
mem[7298] = 80'h0010d7e7c0550102c000;
mem[7299] = 80'h00100001ffabffabffab;
mem[7300] = 80'h0010ff6edf5c0655f137;
mem[7301] = 80'h00101d632caef2926faa;
mem[7302] = 80'h0010b91cd13bf21949e9;
mem[7303] = 80'h01114500000000000000;
mem[7304] = 80'h10100000010000010010;
mem[7305] = 80'h00109400000208004500;
mem[7306] = 80'h0010002f61920000fffd;
mem[7307] = 80'h0010d7e6c0550102c000;
mem[7308] = 80'h00100001ffabffabffab;
mem[7309] = 80'h0010ff6d4d3e733d7b70;
mem[7310] = 80'h0010dd3f5b26c48c1f69;
mem[7311] = 80'h00104bdda96cb2974fd5;
mem[7312] = 80'h0111e300000000000000;
mem[7313] = 80'h00000000000000000000;
mem[7314] = 80'h00000000000000000000;
mem[7315] = 80'h00000000000000000000;
mem[7316] = 80'h10100000010000010010;
mem[7317] = 80'h00109400000208004500;
mem[7318] = 80'h0010002f61930000fffd;
mem[7319] = 80'h0010d7e5c0550102c000;
mem[7320] = 80'h00100001ffabffabffab;
mem[7321] = 80'h0010ff6c3ce05fe502b2;
mem[7322] = 80'h001062f489a12979cf28;
mem[7323] = 80'h00101a929e51c25e63ee;
mem[7324] = 80'h0111fc00000000000000;
mem[7325] = 80'h00000000000000000000;
mem[7326] = 80'h10100000010000010010;
mem[7327] = 80'h00109400000208004500;
mem[7328] = 80'h0010002f61940000fffd;
mem[7329] = 80'h0010d7e4c0550102c000;
mem[7330] = 80'h00100001ffabffabffab;
mem[7331] = 80'h0010ff6b1824b534163d;
mem[7332] = 80'h0010e24c66b045452e6b;
mem[7333] = 80'h0010ff8f5ec10123f185;
mem[7334] = 80'h01111900000000000000;
mem[7335] = 80'h00000000000000000000;
mem[7336] = 80'h00000000000000000000;
mem[7337] = 80'h00000000000000000000;
mem[7338] = 80'h10100000010000010010;
mem[7339] = 80'h00109400000208004500;
mem[7340] = 80'h0010002f61950000fffd;
mem[7341] = 80'h0010d7e3c0550102c000;
mem[7342] = 80'h00100001ffabffabffab;
mem[7343] = 80'h0010ff6a69fa99ec6fff;
mem[7344] = 80'h00105d87b437a8b0feea;
mem[7345] = 80'h0010aed63d7de60bba32;
mem[7346] = 80'h01117d00000000000000;
mem[7347] = 80'h00000000000000000000;
mem[7348] = 80'h10100000010000010010;
mem[7349] = 80'h00109400000208004500;
mem[7350] = 80'h0010002f61960000fffd;
mem[7351] = 80'h0010d7e2c0550102c000;
mem[7352] = 80'h00100001ffabffabffab;
mem[7353] = 80'h0010ff69fb98ec84e5b8;
mem[7354] = 80'h00109ddbc3bf9eae8e69;
mem[7355] = 80'h00105c1a89f1bd28d420;
mem[7356] = 80'h01115600000000000000;
mem[7357] = 80'h00000000000000000000;
mem[7358] = 80'h00000000000000000000;
mem[7359] = 80'h00000000000000000000;
mem[7360] = 80'h00000000000000000000;
mem[7361] = 80'h10100000010000010010;
mem[7362] = 80'h00109400000208004500;
mem[7363] = 80'h0010002f61970000fffd;
mem[7364] = 80'h0010d7e1c0550102c000;
mem[7365] = 80'h00100001ffabffabffab;
mem[7366] = 80'h0010ff688a46c05c9c7a;
mem[7367] = 80'h001022101138735b5e6f;
mem[7368] = 80'h00100dc1e5a520bc3b09;
mem[7369] = 80'h01116300000000000000;
mem[7370] = 80'h10100000010000010010;
mem[7371] = 80'h00109400000208004500;
mem[7372] = 80'h0010002f61980000fffd;
mem[7373] = 80'h0010d7e0c0550102c000;
mem[7374] = 80'h00100001ffabffabffab;
mem[7375] = 80'h0010ff67b2113926cca7;
mem[7376] = 80'h00109caa1d9d46d74c91;
mem[7377] = 80'h001097294fdf1336cf2a;
mem[7378] = 80'h01111d00000000000000;
mem[7379] = 80'h00000000000000000000;
mem[7380] = 80'h00000000000000000000;
mem[7381] = 80'h00000000000000000000;
mem[7382] = 80'h10100000010000010010;
mem[7383] = 80'h00109400000208004500;
mem[7384] = 80'h0010002f61990000fffd;
mem[7385] = 80'h0010d7dfc0550102c000;
mem[7386] = 80'h00100001ffabffabffab;
mem[7387] = 80'h0010ff66c3cf15feb565;
mem[7388] = 80'h00102361cf1aab3d6308;
mem[7389] = 80'h0010c6fadca8cc40ef8b;
mem[7390] = 80'h01111e00000000000000;
mem[7391] = 80'h00000000000000000000;
mem[7392] = 80'h10100000010000010010;
mem[7393] = 80'h00109400000208004500;
mem[7394] = 80'h0010002f619a0000fffd;
mem[7395] = 80'h0010d7dec0550102c000;
mem[7396] = 80'h00100001ffabffabffab;
mem[7397] = 80'h0010ff6551ad60963f22;
mem[7398] = 80'h0010e33db8929d231383;
mem[7399] = 80'h001034bfc1fdcbd9ff15;
mem[7400] = 80'h0111ad00000000000000;
mem[7401] = 80'h00000000000000000000;
mem[7402] = 80'h00000000000000000000;
mem[7403] = 80'h00000000000000000000;
mem[7404] = 80'h10100000010000010010;
mem[7405] = 80'h00109400000208004500;
mem[7406] = 80'h0010002f619b0000fffd;
mem[7407] = 80'h0010d7ddc0550102c000;
mem[7408] = 80'h00100001ffabffabffab;
mem[7409] = 80'h0010ff6420734c4e46e0;
mem[7410] = 80'h00105cf66a1570d6c38a;
mem[7411] = 80'h00106574931858638fe0;
mem[7412] = 80'h01110d00000000000000;
mem[7413] = 80'h00000000000000000000;
mem[7414] = 80'h00000000000000000000;
mem[7415] = 80'h00000000000000000000;
mem[7416] = 80'h10100000010000010010;
mem[7417] = 80'h00109400000208004500;
mem[7418] = 80'h0010002f619c0000fffd;
mem[7419] = 80'h0010d7dcc0550102c000;
mem[7420] = 80'h00100001ffabffabffab;
mem[7421] = 80'h0010ff6304b7a69f526f;
mem[7422] = 80'h0010dc4e85041cea22f1;
mem[7423] = 80'h001080e56fc270d61112;
mem[7424] = 80'h0111b700000000000000;
mem[7425] = 80'h00000000000000000000;
mem[7426] = 80'h10100000010000010010;
mem[7427] = 80'h00109400000208004500;
mem[7428] = 80'h0010002f619d0000fffd;
mem[7429] = 80'h0010d7dbc0550102c000;
mem[7430] = 80'h00100001ffabffabffab;
mem[7431] = 80'h0010ff6275698a472bad;
mem[7432] = 80'h001063855783f11ff288;
mem[7433] = 80'h0010d1266467002df536;
mem[7434] = 80'h01114b00000000000000;
mem[7435] = 80'h00000000000000000000;
mem[7436] = 80'h10100000010000010010;
mem[7437] = 80'h00109400000208004500;
mem[7438] = 80'h0010002f619e0000fffd;
mem[7439] = 80'h0010d7dac0550102c000;
mem[7440] = 80'h00100001ffabffabffab;
mem[7441] = 80'h0010ff61e70bff2fa1ea;
mem[7442] = 80'h0010a3d9200bc70182c2;
mem[7443] = 80'h001023461c892a645502;
mem[7444] = 80'h0111b900000000000000;
mem[7445] = 80'h00000000000000000000;
mem[7446] = 80'h00000000000000000000;
mem[7447] = 80'h00000000000000000000;
mem[7448] = 80'h00000000000000000000;
mem[7449] = 80'h10100000010000010010;
mem[7450] = 80'h00109400000208004500;
mem[7451] = 80'h0010002f619f0000fffd;
mem[7452] = 80'h0010d7d9c0550102c000;
mem[7453] = 80'h00100001ffabffabffab;
mem[7454] = 80'h0010ff6096d5d3f7d828;
mem[7455] = 80'h00101c12f28c2af4528b;
mem[7456] = 80'h00107280820a3cc52305;
mem[7457] = 80'h0111d200000000000000;
mem[7458] = 80'h00000000000000000000;
mem[7459] = 80'h10100000010000010010;
mem[7460] = 80'h00109400000208004500;
mem[7461] = 80'h0010002f61a00000fffd;
mem[7462] = 80'h0010d7d8c0550102c000;
mem[7463] = 80'h00100001ffabffabffab;
mem[7464] = 80'h0010ff5fe5e843761119;
mem[7465] = 80'h001026a6b790cada692a;
mem[7466] = 80'h0010e9525299774296db;
mem[7467] = 80'h01118e00000000000000;
mem[7468] = 80'h00000000000000000000;
mem[7469] = 80'h00000000000000000000;
mem[7470] = 80'h00000000000000000000;
mem[7471] = 80'h10100000010000010010;
mem[7472] = 80'h00109400000208004500;
mem[7473] = 80'h0010002f61a10000fffd;
mem[7474] = 80'h0010d7d7c0550102c000;
mem[7475] = 80'h00100001ffabffabffab;
mem[7476] = 80'h0010ff5e94366fae68db;
mem[7477] = 80'h0010996d6517272fb973;
mem[7478] = 80'h0010b897bf213c57b090;
mem[7479] = 80'h0111c300000000000000;
mem[7480] = 80'h00000000000000000000;
mem[7481] = 80'h10100000010000010010;
mem[7482] = 80'h00109400000208004500;
mem[7483] = 80'h0010002f61a20000fffd;
mem[7484] = 80'h0010d7d6c0550102c000;
mem[7485] = 80'h00100001ffabffabffab;
mem[7486] = 80'h0010ff5d06541ac6e29c;
mem[7487] = 80'h00105931129f1131c838;
mem[7488] = 80'h00104af3c6bda52dcc4e;
mem[7489] = 80'h01119d00000000000000;
mem[7490] = 80'h00000000000000000000;
mem[7491] = 80'h00000000000000000000;
mem[7492] = 80'h00000000000000000000;
mem[7493] = 80'h10100000010000010010;
mem[7494] = 80'h00109400000208004500;
mem[7495] = 80'h0010002f61a30000fffd;
mem[7496] = 80'h0010d7d5c0550102c000;
mem[7497] = 80'h00100001ffabffabffab;
mem[7498] = 80'h0010ff5c778a361e9b5e;
mem[7499] = 80'h0010e6fac018fcc41871;
mem[7500] = 80'h00101b35581d87583954;
mem[7501] = 80'h01116900000000000000;
mem[7502] = 80'h00000000000000000000;
mem[7503] = 80'h10100000010000010010;
mem[7504] = 80'h00109400000208004500;
mem[7505] = 80'h0010002f61a40000fffd;
mem[7506] = 80'h0010d7d4c0550102c000;
mem[7507] = 80'h00100001ffabffabffab;
mem[7508] = 80'h0010ff5b534edccf8fd1;
mem[7509] = 80'h001066422f0990f8f949;
mem[7510] = 80'h0010fefc3b29e6f92061;
mem[7511] = 80'h01116d00000000000000;
mem[7512] = 80'h00000000000000000000;
mem[7513] = 80'h00000000000000000000;
mem[7514] = 80'h00000000000000000000;
mem[7515] = 80'h10100000010000010010;
mem[7516] = 80'h00109400000208004500;
mem[7517] = 80'h0010002f61a50000fffd;
mem[7518] = 80'h0010d7d3c0550102c000;
mem[7519] = 80'h00100001ffabffabffab;
mem[7520] = 80'h0010ff5a2290f017f613;
mem[7521] = 80'h0010d989fd8e7d0d2930;
mem[7522] = 80'h0010af3f30539af95153;
mem[7523] = 80'h01119e00000000000000;
mem[7524] = 80'h00000000000000000000;
mem[7525] = 80'h10100000010000010010;
mem[7526] = 80'h00109400000208004500;
mem[7527] = 80'h0010002f61a60000fffd;
mem[7528] = 80'h0010d7d2c0550102c000;
mem[7529] = 80'h00100001ffabffabffab;
mem[7530] = 80'h0010ff59b0f2857f7c54;
mem[7531] = 80'h001019d58a064b1359bb;
mem[7532] = 80'h00105d7a2dbb79f4b7c1;
mem[7533] = 80'h0111db00000000000000;
mem[7534] = 80'h00000000000000000000;
mem[7535] = 80'h00000000000000000000;
mem[7536] = 80'h00000000000000000000;
mem[7537] = 80'h10100000010000010010;
mem[7538] = 80'h00109400000208004500;
mem[7539] = 80'h0010002f61a70000fffd;
mem[7540] = 80'h0010d7d1c0550102c000;
mem[7541] = 80'h00100001ffabffabffab;
mem[7542] = 80'h0010ff58c12ca9a70596;
mem[7543] = 80'h0010a61e5881a6e68932;
mem[7544] = 80'h00100caae7d96cd9c285;
mem[7545] = 80'h01116100000000000000;
mem[7546] = 80'h00000000000000000000;
mem[7547] = 80'h00000000000000000000;
mem[7548] = 80'h00000000000000000000;
mem[7549] = 80'h10100000010000010010;
mem[7550] = 80'h00109400000208004500;
mem[7551] = 80'h0010002f61a80000fffd;
mem[7552] = 80'h0010d7d0c0550102c000;
mem[7553] = 80'h00100001ffabffabffab;
mem[7554] = 80'h0010ff57f97b50dd554b;
mem[7555] = 80'h001018a45424936a9bcc;
mem[7556] = 80'h001096424dc1e06b91b3;
mem[7557] = 80'h01111300000000000000;
mem[7558] = 80'h10100000010000010010;
mem[7559] = 80'h00109400000208004500;
mem[7560] = 80'h0010002f61a90000fffd;
mem[7561] = 80'h0010d7cfc0550102c000;
mem[7562] = 80'h00100001ffabffabffab;
mem[7563] = 80'h0010ff5688a57c052c89;
mem[7564] = 80'h0010a76f86a37e9f4bd5;
mem[7565] = 80'h0010c78a6c62a2891bd4;
mem[7566] = 80'h01110a00000000000000;
mem[7567] = 80'h00000000000000000000;
mem[7568] = 80'h00000000000000000000;
mem[7569] = 80'h00000000000000000000;
mem[7570] = 80'h10100000010000010010;
mem[7571] = 80'h00109400000208004500;
mem[7572] = 80'h0010002f61aa0000fffd;
mem[7573] = 80'h0010d7cec0550102c000;
mem[7574] = 80'h00100001ffabffabffab;
mem[7575] = 80'h0010ff551ac7096da6ce;
mem[7576] = 80'h00106733f12b48813b5f;
mem[7577] = 80'h001035fc406be236c697;
mem[7578] = 80'h01114b00000000000000;
mem[7579] = 80'h10100000010000010010;
mem[7580] = 80'h00109400000208004500;
mem[7581] = 80'h0010002f61ab0000fffd;
mem[7582] = 80'h0010d7cdc0550102c000;
mem[7583] = 80'h00100001ffabffabffab;
mem[7584] = 80'h0010ff546b1925b5df0c;
mem[7585] = 80'h0010d8f823aca574e8d6;
mem[7586] = 80'h00106475da69c683aca1;
mem[7587] = 80'h01112e00000000000000;
mem[7588] = 80'h00000000000000000000;
mem[7589] = 80'h00000000000000000000;
mem[7590] = 80'h00000000000000000000;
mem[7591] = 80'h10100000010000010010;
mem[7592] = 80'h00109400000208004500;
mem[7593] = 80'h0010002f61ac0000fffd;
mem[7594] = 80'h0010d7ccc0550102c000;
mem[7595] = 80'h00100001ffabffabffab;
mem[7596] = 80'h0010ff534fddcf64cb83;
mem[7597] = 80'h00105840ccbdc94809ad;
mem[7598] = 80'h001081e4260e750fa8e5;
mem[7599] = 80'h0111a200000000000000;
mem[7600] = 80'h00000000000000000000;
mem[7601] = 80'h10100000010000010010;
mem[7602] = 80'h00109400000208004500;
mem[7603] = 80'h0010002f61ad0000fffd;
mem[7604] = 80'h0010d7cbc0550102c000;
mem[7605] = 80'h00100001ffabffabffab;
mem[7606] = 80'h0010ff523e03e3bcb241;
mem[7607] = 80'h0010e78b1e3a24bdd9d4;
mem[7608] = 80'h0010d0272d2c2a217fd2;
mem[7609] = 80'h01118100000000000000;
mem[7610] = 80'h00000000000000000000;
mem[7611] = 80'h00000000000000000000;
mem[7612] = 80'h00000000000000000000;
mem[7613] = 80'h10100000010000010010;
mem[7614] = 80'h00109400000208004500;
mem[7615] = 80'h0010002f61ae0000fffd;
mem[7616] = 80'h0010d7cac0550102c000;
mem[7617] = 80'h00100001ffabffabffab;
mem[7618] = 80'h0010ff51ac6196d43806;
mem[7619] = 80'h001027d769b212a3a91f;
mem[7620] = 80'h0010226ffcb6188fdd1a;
mem[7621] = 80'h01114d00000000000000;
mem[7622] = 80'h00000000000000000000;
mem[7623] = 80'h10100000010000010010;
mem[7624] = 80'h00109400000208004500;
mem[7625] = 80'h0010002f61af0000fffd;
mem[7626] = 80'h0010d7c9c0550102c000;
mem[7627] = 80'h00100001ffabffabffab;
mem[7628] = 80'h0010ff50ddbfba0c41c4;
mem[7629] = 80'h0010981cbb35ff567956;
mem[7630] = 80'h001073a9627584158e09;
mem[7631] = 80'h0111db00000000000000;
mem[7632] = 80'h00000000000000000000;
mem[7633] = 80'h00000000000000000000;
mem[7634] = 80'h00000000000000000000;
mem[7635] = 80'h10100000010000010010;
mem[7636] = 80'h00109400000208004500;
mem[7637] = 80'h0010002f61b00000fffd;
mem[7638] = 80'h0010d7c8c0550102c000;
mem[7639] = 80'h00100001ffabffabffab;
mem[7640] = 80'h0010ff4fdcce642099bd;
mem[7641] = 80'h00105aa370f879bb8c65;
mem[7642] = 80'h0010162c861ab7940f26;
mem[7643] = 80'h01111700000000000000;
mem[7644] = 80'h00000000000000000000;
mem[7645] = 80'h10100000010000010010;
mem[7646] = 80'h00109400000208004500;
mem[7647] = 80'h0010002f61b10000fffd;
mem[7648] = 80'h0010d7c7c0550102c000;
mem[7649] = 80'h00100001ffabffabffab;
mem[7650] = 80'h0010ff4ead1048f8e07f;
mem[7651] = 80'h0010e568a27f944e5c24;
mem[7652] = 80'h00104763b169b8c2c4ad;
mem[7653] = 80'h0111ee00000000000000;
mem[7654] = 80'h00000000000000000000;
mem[7655] = 80'h00000000000000000000;
mem[7656] = 80'h00000000000000000000;
mem[7657] = 80'h10100000010000010010;
mem[7658] = 80'h00109400000208004500;
mem[7659] = 80'h0010002f61b20000fffd;
mem[7660] = 80'h0010d7c6c0550102c000;
mem[7661] = 80'h00100001ffabffabffab;
mem[7662] = 80'h0010ff4d3f723d906a38;
mem[7663] = 80'h00102534d5f7a2502cf7;
mem[7664] = 80'h0010b5a1ba61de567d6b;
mem[7665] = 80'h0111e000000000000000;
mem[7666] = 80'h00000000000000000000;
mem[7667] = 80'h10100000010000010010;
mem[7668] = 80'h00109400000208004500;
mem[7669] = 80'h0010002f61b30000fffd;
mem[7670] = 80'h0010d7c5c0550102c000;
mem[7671] = 80'h00100001ffabffabffab;
mem[7672] = 80'h0010ff4c4eac114813fa;
mem[7673] = 80'h00109aff07704fa5fcb6;
mem[7674] = 80'h0010e4ee8d0a2be2dc63;
mem[7675] = 80'h01118e00000000000000;
mem[7676] = 80'h00000000000000000000;
mem[7677] = 80'h00000000000000000000;
mem[7678] = 80'h00000000000000000000;
mem[7679] = 80'h10100000010000010010;
mem[7680] = 80'h00109400000208004500;
mem[7681] = 80'h0010002f61b40000fffd;
mem[7682] = 80'h0010d7c4c0550102c000;
mem[7683] = 80'h00100001ffabffabffab;
mem[7684] = 80'h0010ff4b6a68fb990775;
mem[7685] = 80'h00101a47e86123991c05;
mem[7686] = 80'h001001d7bc1e92d1b884;
mem[7687] = 80'h0111ac00000000000000;
mem[7688] = 80'h00000000000000000000;
mem[7689] = 80'h10100000010000010010;
mem[7690] = 80'h00109400000208004500;
mem[7691] = 80'h0010002f61b50000fffd;
mem[7692] = 80'h0010d7c3c0550102c000;
mem[7693] = 80'h00100001ffabffabffab;
mem[7694] = 80'h0010ff4a1bb6d7417eb7;
mem[7695] = 80'h0010a58c3ae6ce6ccc44;
mem[7696] = 80'h001050988b4937f96944;
mem[7697] = 80'h0111e200000000000000;
mem[7698] = 80'h00000000000000000000;
mem[7699] = 80'h00000000000000000000;
mem[7700] = 80'h00000000000000000000;
mem[7701] = 80'h00000000000000000000;
mem[7702] = 80'h10100000010000010010;
mem[7703] = 80'h00109400000208004500;
mem[7704] = 80'h0010002f61b60000fffd;
mem[7705] = 80'h0010d7c2c0550102c000;
mem[7706] = 80'h00100001ffabffabffab;
mem[7707] = 80'h0010ff4989d4a229f4f0;
mem[7708] = 80'h001065d04d6ef872bcf7;
mem[7709] = 80'h0010a251aacc2908845e;
mem[7710] = 80'h0111d600000000000000;
mem[7711] = 80'h00000000000000000000;
mem[7712] = 80'h10100000010000010010;
mem[7713] = 80'h00109400000208004500;
mem[7714] = 80'h0010002f61b70000fffd;
mem[7715] = 80'h0010d7c1c0550102c000;
mem[7716] = 80'h00100001ffabffabffab;
mem[7717] = 80'h0010ff48f80a8ef18d32;
mem[7718] = 80'h0010da1b9fe915876cf7;
mem[7719] = 80'h0010f32060e39b56cd17;
mem[7720] = 80'h0111ad00000000000000;
mem[7721] = 80'h00000000000000000000;
mem[7722] = 80'h00000000000000000000;
mem[7723] = 80'h00000000000000000000;
mem[7724] = 80'h10100000010000010010;
mem[7725] = 80'h00109400000208004500;
mem[7726] = 80'h0010002f61b80000fffd;
mem[7727] = 80'h0010d7c0c0550102c000;
mem[7728] = 80'h00100001ffabffabffab;
mem[7729] = 80'h0010ff47c05d778bddef;
mem[7730] = 80'h001064a1934c200b7e01;
mem[7731] = 80'h0010694163a387cfc7e7;
mem[7732] = 80'h0111f700000000000000;
mem[7733] = 80'h00000000000000000000;
mem[7734] = 80'h10100000010000010010;
mem[7735] = 80'h00109400000208004500;
mem[7736] = 80'h0010002f61b90000fffd;
mem[7737] = 80'h0010d7bfc0550102c000;
mem[7738] = 80'h00100001ffabffabffab;
mem[7739] = 80'h0010ff46b1835b53a42d;
mem[7740] = 80'h0010db6a41cbcdfeae80;
mem[7741] = 80'h0010381800e77c642fc1;
mem[7742] = 80'h0111e000000000000000;
mem[7743] = 80'h00000000000000000000;
mem[7744] = 80'h00000000000000000000;
mem[7745] = 80'h00000000000000000000;
mem[7746] = 80'h10100000010000010010;
mem[7747] = 80'h00109400000208004500;
mem[7748] = 80'h0010002f61ba0000fffd;
mem[7749] = 80'h0010d7bec0550102c000;
mem[7750] = 80'h00100001ffabffabffab;
mem[7751] = 80'h0010ff4523e12e3b2e6a;
mem[7752] = 80'h00101b363643fbe0de13;
mem[7753] = 80'h0010cad7c7edc1bb42b7;
mem[7754] = 80'h0111a800000000000000;
mem[7755] = 80'h00000000000000000000;
mem[7756] = 80'h10100000010000010010;
mem[7757] = 80'h00109400000208004500;
mem[7758] = 80'h0010002f61bb0000fffd;
mem[7759] = 80'h0010d7bdc0550102c000;
mem[7760] = 80'h00100001ffabffabffab;
mem[7761] = 80'h0010ff44523f02e357a8;
mem[7762] = 80'h0010a4fde4c416150e12;
mem[7763] = 80'h00109b953c71cd5863a4;
mem[7764] = 80'h01113c00000000000000;
mem[7765] = 80'h00000000000000000000;
mem[7766] = 80'h00000000000000000000;
mem[7767] = 80'h00000000000000000000;
mem[7768] = 80'h10100000010000010010;
mem[7769] = 80'h00109400000208004500;
mem[7770] = 80'h0010002f61bc0000fffd;
mem[7771] = 80'h0010d7bcc0550102c000;
mem[7772] = 80'h00100001ffabffabffab;
mem[7773] = 80'h0010ff4376fbe8324327;
mem[7774] = 80'h001024450bd57a29ef61;
mem[7775] = 80'h00107e8d6933dcc46860;
mem[7776] = 80'h0111ca00000000000000;
mem[7777] = 80'h00000000000000000000;
mem[7778] = 80'h10100000010000010010;
mem[7779] = 80'h00109400000208004500;
mem[7780] = 80'h0010002f61bd0000fffd;
mem[7781] = 80'h0010d7bbc0550102c000;
mem[7782] = 80'h00100001ffabffabffab;
mem[7783] = 80'h0010ff420725c4ea3ae5;
mem[7784] = 80'h00109b8ed95297dc38e3;
mem[7785] = 80'h00102f04c922bbc8bf48;
mem[7786] = 80'h0111ae00000000000000;
mem[7787] = 80'h00000000000000000000;
mem[7788] = 80'h00000000000000000000;
mem[7789] = 80'h00000000000000000000;
mem[7790] = 80'h10100000010000010010;
mem[7791] = 80'h00109400000208004500;
mem[7792] = 80'h0010002f61be0000fffd;
mem[7793] = 80'h0010d7bac0550102c000;
mem[7794] = 80'h00100001ffabffabffab;
mem[7795] = 80'h0010ff419547b182b0a2;
mem[7796] = 80'h00105bd2aedaa1c24850;
mem[7797] = 80'h0010ddcde8c34dd09612;
mem[7798] = 80'h01113500000000000000;
mem[7799] = 80'h00000000000000000000;
mem[7800] = 80'h10100000010000010010;
mem[7801] = 80'h00109400000208004500;
mem[7802] = 80'h0010002f61bf0000fffd;
mem[7803] = 80'h0010d7b9c0550102c000;
mem[7804] = 80'h00100001ffabffabffab;
mem[7805] = 80'h0010ff40e4999d5ac960;
mem[7806] = 80'h0010e4197c5d4c379811;
mem[7807] = 80'h00108c82df2704474cd6;
mem[7808] = 80'h01112500000000000000;
mem[7809] = 80'h00000000000000000000;
mem[7810] = 80'h00000000000000000000;
mem[7811] = 80'h00000000000000000000;
mem[7812] = 80'h10100000010000010010;
mem[7813] = 80'h00109400000208004500;
mem[7814] = 80'h0010002f61c00000fffd;
mem[7815] = 80'h0010d7b8c0550102c000;
mem[7816] = 80'h00100001ffabffabffab;
mem[7817] = 80'h0010ff3f733c908122c0;
mem[7818] = 80'h00102eba24e3619e3f93;
mem[7819] = 80'h0010eb63f10f0808833f;
mem[7820] = 80'h01117800000000000000;
mem[7821] = 80'h00000000000000000000;
mem[7822] = 80'h10100000010000010010;
mem[7823] = 80'h00109400000208004500;
mem[7824] = 80'h0010002f61c10000fffd;
mem[7825] = 80'h0010d7b7c0550102c000;
mem[7826] = 80'h00100001ffabffabffab;
mem[7827] = 80'h0010ff3e02e2bc595b02;
mem[7828] = 80'h00109171f6648c6befd2;
mem[7829] = 80'h0010ba2cc641618dc48d;
mem[7830] = 80'h01114f00000000000000;
mem[7831] = 80'h00000000000000000000;
mem[7832] = 80'h00000000000000000000;
mem[7833] = 80'h00000000000000000000;
mem[7834] = 80'h10100000010000010010;
mem[7835] = 80'h00109400000208004500;
mem[7836] = 80'h0010002f61c20000fffd;
mem[7837] = 80'h0010d7b6c0550102c000;
mem[7838] = 80'h00100001ffabffabffab;
mem[7839] = 80'h0010ff3d9080c931d145;
mem[7840] = 80'h0010512d81ecba759f81;
mem[7841] = 80'h001048f555c409169b76;
mem[7842] = 80'h01114200000000000000;
mem[7843] = 80'h00000000000000000000;
mem[7844] = 80'h10100000010000010010;
mem[7845] = 80'h00109400000208004500;
mem[7846] = 80'h0010002f61c30000fffd;
mem[7847] = 80'h0010d7b5c0550102c000;
mem[7848] = 80'h00100001ffabffabffab;
mem[7849] = 80'h0010ff3ce15ee5e9a887;
mem[7850] = 80'h0010eee6536b57804fc1;
mem[7851] = 80'h0010198953d6396fc5e6;
mem[7852] = 80'h01113500000000000000;
mem[7853] = 80'h00000000000000000000;
mem[7854] = 80'h00000000000000000000;
mem[7855] = 80'h00000000000000000000;
mem[7856] = 80'h10100000010000010010;
mem[7857] = 80'h00109400000208004500;
mem[7858] = 80'h0010002f61c40000fffd;
mem[7859] = 80'h0010d7b4c0550102c000;
mem[7860] = 80'h00100001ffabffabffab;
mem[7861] = 80'h0010ff3bc59a0f38bc08;
mem[7862] = 80'h00106e5ebc7a3bbcaef2;
mem[7863] = 80'h0010fc9ccac39267e2eb;
mem[7864] = 80'h01117800000000000000;
mem[7865] = 80'h00000000000000000000;
mem[7866] = 80'h10100000010000010010;
mem[7867] = 80'h00109400000208004500;
mem[7868] = 80'h0010002f61c50000fffd;
mem[7869] = 80'h0010d7b3c0550102c000;
mem[7870] = 80'h00100001ffabffabffab;
mem[7871] = 80'h0010ff3ab44423e0c5ca;
mem[7872] = 80'h0010d1956efdd6497eb3;
mem[7873] = 80'h0010add3fd7121b781f6;
mem[7874] = 80'h0111e100000000000000;
mem[7875] = 80'h00000000000000000000;
mem[7876] = 80'h00000000000000000000;
mem[7877] = 80'h00000000000000000000;
mem[7878] = 80'h10100000010000010010;
mem[7879] = 80'h00109400000208004500;
mem[7880] = 80'h0010002f61c60000fffd;
mem[7881] = 80'h0010d7b2c0550102c000;
mem[7882] = 80'h00100001ffabffabffab;
mem[7883] = 80'h0010ff39262656884f8d;
mem[7884] = 80'h001011c91975e0570e00;
mem[7885] = 80'h00105f1adcd9de47e4cb;
mem[7886] = 80'h01112200000000000000;
mem[7887] = 80'h00000000000000000000;
mem[7888] = 80'h10100000010000010010;
mem[7889] = 80'h00109400000208004500;
mem[7890] = 80'h0010002f61c70000fffd;
mem[7891] = 80'h0010d7b1c0550102c000;
mem[7892] = 80'h00100001ffabffabffab;
mem[7893] = 80'h0010ff3857f87a50364f;
mem[7894] = 80'h0010ae02cbf20da2df81;
mem[7895] = 80'h00100e748fa1f2b6d0ec;
mem[7896] = 80'h01113200000000000000;
mem[7897] = 80'h00000000000000000000;
mem[7898] = 80'h00000000000000000000;
mem[7899] = 80'h00000000000000000000;
mem[7900] = 80'h10100000010000010010;
mem[7901] = 80'h00109400000208004500;
mem[7902] = 80'h0010002f61c80000fffd;
mem[7903] = 80'h0010d7b0c0550102c000;
mem[7904] = 80'h00100001ffabffabffab;
mem[7905] = 80'h0010ff376faf832a6692;
mem[7906] = 80'h001010b8c757382ecd77;
mem[7907] = 80'h001094158c90a83d7687;
mem[7908] = 80'h0111c100000000000000;
mem[7909] = 80'h10100000010000010010;
mem[7910] = 80'h00109400000208004500;
mem[7911] = 80'h0010002f61c90000fffd;
mem[7912] = 80'h0010d7afc0550102c000;
mem[7913] = 80'h00100001ffabffabffab;
mem[7914] = 80'h0010ff361e71aff21f50;
mem[7915] = 80'h0010af7315d0d5db1d71;
mem[7916] = 80'h0010c5cee0b5b3ee7ce0;
mem[7917] = 80'h01116f00000000000000;
mem[7918] = 80'h00000000000000000000;
mem[7919] = 80'h00000000000000000000;
mem[7920] = 80'h00000000000000000000;
mem[7921] = 80'h10100000010000010010;
mem[7922] = 80'h00109400000208004500;
mem[7923] = 80'h0010002f61ca0000fffd;
mem[7924] = 80'h0010d7aec0550102c000;
mem[7925] = 80'h00100001ffabffabffab;
mem[7926] = 80'h0010ff358c13da9a9517;
mem[7927] = 80'h00106f2f6258e3c56dfa;
mem[7928] = 80'h0010378bfd30ac3e312a;
mem[7929] = 80'h01114e00000000000000;
mem[7930] = 80'h00000000000000000000;
mem[7931] = 80'h00000000000000000000;
mem[7932] = 80'h00000000000000000000;
mem[7933] = 80'h10100000010000010010;
mem[7934] = 80'h00109400000208004500;
mem[7935] = 80'h0010002f61cb0000fffd;
mem[7936] = 80'h0010d7adc0550102c000;
mem[7937] = 80'h00100001ffabffabffab;
mem[7938] = 80'h0010ff34fdcdf642ecd5;
mem[7939] = 80'h0010d0e4b0df0e30bd63;
mem[7940] = 80'h001066584434270d4daa;
mem[7941] = 80'h01119700000000000000;
mem[7942] = 80'h10100000010000010010;
mem[7943] = 80'h00109400000208004500;
mem[7944] = 80'h0010002f61cc0000fffd;
mem[7945] = 80'h0010d7acc0550102c000;
mem[7946] = 80'h00100001ffabffabffab;
mem[7947] = 80'h0010ff33d9091c93f85a;
mem[7948] = 80'h0010505c5fce620c5c18;
mem[7949] = 80'h001083c9b8bb67c393fd;
mem[7950] = 80'h0111a900000000000000;
mem[7951] = 80'h00000000000000000000;
mem[7952] = 80'h00000000000000000000;
mem[7953] = 80'h00000000000000000000;
mem[7954] = 80'h10100000010000010010;
mem[7955] = 80'h00109400000208004500;
mem[7956] = 80'h0010002f61cd0000fffd;
mem[7957] = 80'h0010d7abc0550102c000;
mem[7958] = 80'h00100001ffabffabffab;
mem[7959] = 80'h0010ff32a8d7304b8198;
mem[7960] = 80'h0010ef978d498ff98c11;
mem[7961] = 80'h0010d202ea2250e5ea69;
mem[7962] = 80'h01116300000000000000;
mem[7963] = 80'h00000000000000000000;
mem[7964] = 80'h10100000010000010010;
mem[7965] = 80'h00109400000208004500;
mem[7966] = 80'h0010002f61ce0000fffd;
mem[7967] = 80'h0010d7aac0550102c000;
mem[7968] = 80'h00100001ffabffabffab;
mem[7969] = 80'h0010ff313ab545230bdf;
mem[7970] = 80'h00102fcbfac1b9e7fc9a;
mem[7971] = 80'h00102047f7bf7bd9cb0c;
mem[7972] = 80'h0111e100000000000000;
mem[7973] = 80'h00000000000000000000;
mem[7974] = 80'h00000000000000000000;
mem[7975] = 80'h00000000000000000000;
mem[7976] = 80'h10100000010000010010;
mem[7977] = 80'h00109400000208004500;
mem[7978] = 80'h0010002f61cf0000fffd;
mem[7979] = 80'h0010d7a9c0550102c000;
mem[7980] = 80'h00100001ffabffabffab;
mem[7981] = 80'h0010ff304b6b69fb721d;
mem[7982] = 80'h00109000284654122ce3;
mem[7983] = 80'h00107184fc8a311d2435;
mem[7984] = 80'h01119200000000000000;
mem[7985] = 80'h00000000000000000000;
mem[7986] = 80'h10100000010000010010;
mem[7987] = 80'h00109400000208004500;
mem[7988] = 80'h0010002f61d00000fffd;
mem[7989] = 80'h0010d7a8c0550102c000;
mem[7990] = 80'h00100001ffabffabffab;
mem[7991] = 80'h0010ff2f4a1ab7d7aa64;
mem[7992] = 80'h001052bfe38bd2ffdad6;
mem[7993] = 80'h001014f2ee656c233eb8;
mem[7994] = 80'h01110d00000000000000;
mem[7995] = 80'h00000000000000000000;
mem[7996] = 80'h00000000000000000000;
mem[7997] = 80'h00000000000000000000;
mem[7998] = 80'h00000000000000000000;
mem[7999] = 80'h10100000010000010010;
mem[8000] = 80'h00109400000208004500;
mem[8001] = 80'h0010002f61d10000fffd;
mem[8002] = 80'h0010d7a7c0550102c000;
mem[8003] = 80'h00100001ffabffabffab;
mem[8004] = 80'h0010ff2e3bc49b0fd3a6;
mem[8005] = 80'h0010ed74310c3f0a0a9f;
mem[8006] = 80'h0010453470f837c9a363;
mem[8007] = 80'h0111f200000000000000;
mem[8008] = 80'h10100000010000010010;
mem[8009] = 80'h00109400000208004500;
mem[8010] = 80'h0010002f61d20000fffd;
mem[8011] = 80'h0010d7a6c0550102c000;
mem[8012] = 80'h00100001ffabffabffab;
mem[8013] = 80'h0010ff2da9a6ee6759e1;
mem[8014] = 80'h00102d28468409147a54;
mem[8015] = 80'h0010b77ca150be123f68;
mem[8016] = 80'h01118f00000000000000;
mem[8017] = 80'h00000000000000000000;
mem[8018] = 80'h00000000000000000000;
mem[8019] = 80'h00000000000000000000;
mem[8020] = 80'h10100000010000010010;
mem[8021] = 80'h00109400000208004500;
mem[8022] = 80'h0010002f61d30000fffd;
mem[8023] = 80'h0010d7a5c0550102c000;
mem[8024] = 80'h00100001ffabffabffab;
mem[8025] = 80'h0010ff2cd878c2bf2023;
mem[8026] = 80'h001092e39403e4e1aa0d;
mem[8027] = 80'h0010e6b94ce75b9e6225;
mem[8028] = 80'h01113c00000000000000;
mem[8029] = 80'h00000000000000000000;
mem[8030] = 80'h10100000010000010010;
mem[8031] = 80'h00109400000208004500;
mem[8032] = 80'h0010002f61d40000fffd;
mem[8033] = 80'h0010d7a4c0550102c000;
mem[8034] = 80'h00100001ffabffabffab;
mem[8035] = 80'h0010ff2bfcbc286e34ac;
mem[8036] = 80'h0010125b7b1288dd4bb6;
mem[8037] = 80'h0010033ee4bd5ca2c9aa;
mem[8038] = 80'h01111900000000000000;
mem[8039] = 80'h00000000000000000000;
mem[8040] = 80'h00000000000000000000;
mem[8041] = 80'h00000000000000000000;
mem[8042] = 80'h10100000010000010010;
mem[8043] = 80'h00109400000208004500;
mem[8044] = 80'h0010002f61d50000fffd;
mem[8045] = 80'h0010d7a3c0550102c000;
mem[8046] = 80'h00100001ffabffabffab;
mem[8047] = 80'h0010ff2a8d6204b64d6e;
mem[8048] = 80'h0010ad90a99565289bff;
mem[8049] = 80'h001052f87a07fb34e91f;
mem[8050] = 80'h0111f800000000000000;
mem[8051] = 80'h00000000000000000000;
mem[8052] = 80'h10100000010000010010;
mem[8053] = 80'h00109400000208004500;
mem[8054] = 80'h0010002f61d60000fffd;
mem[8055] = 80'h0010d7a2c0550102c000;
mem[8056] = 80'h00100001ffabffabffab;
mem[8057] = 80'h0010ff291f0071dec729;
mem[8058] = 80'h00106dccde1d5336eb37;
mem[8059] = 80'h0010a0e5f88f84b31bf3;
mem[8060] = 80'h01115000000000000000;
mem[8061] = 80'h00000000000000000000;
mem[8062] = 80'h00000000000000000000;
mem[8063] = 80'h00000000000000000000;
mem[8064] = 80'h00000000000000000000;
mem[8065] = 80'h10100000010000010010;
mem[8066] = 80'h00109400000208004500;
mem[8067] = 80'h0010002f61d70000fffd;
mem[8068] = 80'h0010d7a1c0550102c000;
mem[8069] = 80'h00100001ffabffabffab;
mem[8070] = 80'h0010ff286ede5d06beeb;
mem[8071] = 80'h0010d2070c9abec33b4e;
mem[8072] = 80'h0010f126f32bb8259bf6;
mem[8073] = 80'h0111f200000000000000;
mem[8074] = 80'h10100000010000010010;
mem[8075] = 80'h00109400000208004500;
mem[8076] = 80'h0010002f61d80000fffd;
mem[8077] = 80'h0010d7a0c0550102c000;
mem[8078] = 80'h00100001ffabffabffab;
mem[8079] = 80'h0010ff275689a47cee36;
mem[8080] = 80'h00106cbd003f8b4f29b0;
mem[8081] = 80'h00106bce59d12f1590ed;
mem[8082] = 80'h01116600000000000000;
mem[8083] = 80'h00000000000000000000;
mem[8084] = 80'h00000000000000000000;
mem[8085] = 80'h00000000000000000000;
mem[8086] = 80'h10100000010000010010;
mem[8087] = 80'h00109400000208004500;
mem[8088] = 80'h0010002f61d90000fffd;
mem[8089] = 80'h0010d79fc0550102c000;
mem[8090] = 80'h00100001ffabffabffab;
mem[8091] = 80'h0010ff26275788a497f4;
mem[8092] = 80'h0010d376d2b866baf839;
mem[8093] = 80'h00103a29a39bd55bd3e3;
mem[8094] = 80'h0111ee00000000000000;
mem[8095] = 80'h00000000000000000000;
mem[8096] = 80'h10100000010000010010;
mem[8097] = 80'h00109400000208004500;
mem[8098] = 80'h0010002f61da0000fffd;
mem[8099] = 80'h0010d79ec0550102c000;
mem[8100] = 80'h00100001ffabffabffab;
mem[8101] = 80'h0010ff25b535fdcc1db3;
mem[8102] = 80'h0010132aa53050a488b2;
mem[8103] = 80'h0010c86cbe0617bba850;
mem[8104] = 80'h0111b500000000000000;
mem[8105] = 80'h00000000000000000000;
mem[8106] = 80'h00000000000000000000;
mem[8107] = 80'h00000000000000000000;
mem[8108] = 80'h10100000010000010010;
mem[8109] = 80'h00109400000208004500;
mem[8110] = 80'h0010002f61db0000fffd;
mem[8111] = 80'h0010d79dc0550102c000;
mem[8112] = 80'h00100001ffabffabffab;
mem[8113] = 80'h0010ff24c4ebd1146471;
mem[8114] = 80'h0010ace177b7bd5158ab;
mem[8115] = 80'h001099a49f2e922fbff1;
mem[8116] = 80'h0111d800000000000000;
mem[8117] = 80'h00000000000000000000;
mem[8118] = 80'h00000000000000000000;
mem[8119] = 80'h00000000000000000000;
mem[8120] = 80'h10100000010000010010;
mem[8121] = 80'h00109400000208004500;
mem[8122] = 80'h0010002f61dc0000fffd;
mem[8123] = 80'h0010d79cc0550102c000;
mem[8124] = 80'h00100001ffabffabffab;
mem[8125] = 80'h0010ff23e02f3bc570fe;
mem[8126] = 80'h00102c5998a6d16db9d1;
mem[8127] = 80'h00107c0652a3543b2e20;
mem[8128] = 80'h0111dc00000000000000;
mem[8129] = 80'h00000000000000000000;
mem[8130] = 80'h10100000010000010010;
mem[8131] = 80'h00109400000208004500;
mem[8132] = 80'h0010002f61dd0000fffd;
mem[8133] = 80'h0010d79bc0550102c000;
mem[8134] = 80'h00100001ffabffabffab;
mem[8135] = 80'h0010ff2291f1171d093c;
mem[8136] = 80'h001093924a213c986958;
mem[8137] = 80'h00102dd6981804c8c878;
mem[8138] = 80'h01110800000000000000;
mem[8139] = 80'h00000000000000000000;
mem[8140] = 80'h10100000010000010010;
mem[8141] = 80'h00109400000208004500;
mem[8142] = 80'h0010002f61de0000fffd;
mem[8143] = 80'h0010d79ac0550102c000;
mem[8144] = 80'h00100001ffabffabffab;
mem[8145] = 80'h0010ff2103936275837b;
mem[8146] = 80'h001053ce3da90a8619d3;
mem[8147] = 80'h0010df9385f5fbcf869c;
mem[8148] = 80'h01112400000000000000;
mem[8149] = 80'h00000000000000000000;
mem[8150] = 80'h00000000000000000000;
mem[8151] = 80'h00000000000000000000;
mem[8152] = 80'h00000000000000000000;
mem[8153] = 80'h10100000010000010010;
mem[8154] = 80'h00109400000208004500;
mem[8155] = 80'h0010002f61df0000fffd;
mem[8156] = 80'h0010d799c0550102c000;
mem[8157] = 80'h00100001ffabffabffab;
mem[8158] = 80'h0010ff20724d4eadfab9;
mem[8159] = 80'h0010ec05ef2ee773c9aa;
mem[8160] = 80'h00108e508e869b5e483d;
mem[8161] = 80'h01112a00000000000000;
mem[8162] = 80'h00000000000000000000;
mem[8163] = 80'h10100000010000010010;
mem[8164] = 80'h00109400000208004500;
mem[8165] = 80'h0010002f61e00000fffd;
mem[8166] = 80'h0010d798c0550102c000;
mem[8167] = 80'h00100001ffabffabffab;
mem[8168] = 80'h0010ff1f0170de2c3388;
mem[8169] = 80'h0010d6b1aa32075df20b;
mem[8170] = 80'h001015825eebfe253c0a;
mem[8171] = 80'h01112000000000000000;
mem[8172] = 80'h00000000000000000000;
mem[8173] = 80'h00000000000000000000;
mem[8174] = 80'h00000000000000000000;
mem[8175] = 80'h10100000010000010010;
mem[8176] = 80'h00109400000208004500;
mem[8177] = 80'h0010002f61e10000fffd;
mem[8178] = 80'h0010d797c0550102c000;
mem[8179] = 80'h00100001ffabffabffab;
mem[8180] = 80'h0010ff1e70aef2f44a4a;
mem[8181] = 80'h0010697a78b5eaa82242;
mem[8182] = 80'h00104444c0945e351bf6;
mem[8183] = 80'h01119900000000000000;
mem[8184] = 80'h00000000000000000000;
mem[8185] = 80'h00000000000000000000;
mem[8186] = 80'h00000000000000000000;
mem[8187] = 80'h00000000000000000000;
mem[8188] = 80'h00000000000000000000;
mem[8189] = 80'h00000000000000000000;
mem[8190] = 80'h00000000000000000000;
mem[8191] = 80'h00000000000000000000;
end


//*********************
//MAIN CORE
//********************* 
reg [15:0] time_cnt ;    
reg [31:0] cnt ;

initial begin
    time_cnt = 'd0 ;
    cnt      = 'd0 ;
end

always @(posedge clk) begin

    if ( time_cnt == 'd1000 ) begin
        time_cnt <= time_cnt ;
    end
    else begin
        time_cnt <= time_cnt+1'b1 ;
    end
end

always @(posedge clk) begin

    if ( time_cnt >'d900 ) begin
        if ( cnt == 'd8191 ) begin
            cnt <= 'd0 ;
        end
        else begin
           cnt <= cnt+1'b1 ; 
        end
    end
    else begin
        cnt <= 'd0 ;
    end
end

wire [12:0] rd_addr ;

assign rd_addr = cnt[12:0] ;


always @(posedge clk) begin
	dout_ff <= mem[rd_addr] ;
end


assign sop  = dout_ff[76] ;
assign eop  = dout_ff[72] ;
assign dval = dout_ff[68] ;
assign mod  = dout_ff[66:64] ;
assign dout = dout_ff[63:0] ;


//*********************
endmodule   